module uncache (
    input 
);
    
endmodule