module uncache (

);
    
endmodule