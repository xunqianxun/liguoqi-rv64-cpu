/************************************************************
Author:LiGuoqi
Name:mmio.v
Function:memory mapped I/O
************************************************************/
module mmio (
    input         wire                                  clk             ,
    input         wire                                  rst             ,

    
);
    
endmodule