module top(
  input wire a,
  input wire b,
  output wire  f
);
  assign f = a ^ b;
endmodule
