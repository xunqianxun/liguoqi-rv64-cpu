/************************************************************
Author:LiGuoqi
Name:arbitrate.v
Function:arbitrate i_cache and d_cache
************************************************************/
module arbitrate (
    input       wire                                         clk            ,
    input       wire                                         rst            ,

    
);
    
endmodule