/* verilator lint_off DECLFILENAME */
/* verilator lint_off UNUSED */
module ysyx_210340_InstFetch(
  input         clock,
  input         reset,
  input         io_stall,
  input         io_flush,
  input         io_br_en,
  input  [31:0] io_br_addr,
  output [31:0] io_out_pc,
  output [31:0] io_out_inst,
  output        io_out_imem_hs,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output [31:0] io_imem_req_bits_addr,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[InstFetch.scala 19:22]
  reg [31:0] pc; // @[InstFetch.scala 25:19]
  wire [31:0] _pc_nxt_T_1 = pc + 32'h4; // @[InstFetch.scala 26:45]
  wire [31:0] pc_nxt = io_br_en ? io_br_addr : _pc_nxt_T_1; // @[InstFetch.scala 26:19]
  reg [31:0] inst; // @[InstFetch.scala 27:21]
  wire  _io_imem_req_valid_T_1 = ~io_stall; // @[InstFetch.scala 36:37]
  wire  _T = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_2 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _state_T_2 = io_flush ? 2'h1 : 2'h3; // @[InstFetch.scala 54:19]
  wire [1:0] _GEN_0 = _io_imem_req_valid_T_1 & _T_4 ? _state_T_2 : state; // @[InstFetch.scala 52:35 InstFetch.scala 54:13 InstFetch.scala 19:22]
  wire  _T_6 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_7 = io_imem_resp_ready & io_imem_resp_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _inst_T_6 = pc[2] ? io_imem_resp_bits_rdata[63:32] : io_imem_resp_bits_rdata[31:0]; // @[InstFetch.scala 61:75]
  wire [31:0] _inst_T_7 = ~io_imem_req_bits_addr[31] ? io_imem_resp_bits_rdata[31:0] : _inst_T_6; // @[InstFetch.scala 61:20]
  wire [31:0] _GEN_1 = _T_7 ? _inst_T_7 : inst; // @[InstFetch.scala 59:26 InstFetch.scala 61:14 InstFetch.scala 27:21]
  wire [1:0] _GEN_2 = _T_7 ? 2'h1 : _state_T_2; // @[InstFetch.scala 59:26 InstFetch.scala 63:17 InstFetch.scala 58:13]
  wire [1:0] _GEN_3 = _T_6 ? _GEN_2 : state; // @[Conditional.scala 39:67 InstFetch.scala 19:22]
  wire [31:0] _GEN_4 = _T_6 ? _GEN_1 : inst; // @[Conditional.scala 39:67 InstFetch.scala 27:21]
  wire  _io_out_pc_T = state == 2'h1; // @[InstFetch.scala 68:27]
  reg  io_out_pc_REG; // @[InstFetch.scala 68:49]
  reg  io_out_inst_REG; // @[InstFetch.scala 69:51]
  assign io_out_pc = state == 2'h1 & io_out_pc_REG ? pc : 32'h0; // @[InstFetch.scala 68:19]
  assign io_out_inst = _io_out_pc_T & io_out_inst_REG ? inst : 32'h0; // @[InstFetch.scala 69:21]
  assign io_out_imem_hs = io_imem_resp_valid & io_imem_resp_ready; // @[InstFetch.scala 70:32]
  assign io_imem_req_valid = state == 2'h2 & ~io_stall; // @[InstFetch.scala 36:34]
  assign io_imem_req_bits_addr = pc; // @[InstFetch.scala 30:17]
  assign io_imem_resp_ready = state == 2'h3; // @[InstFetch.scala 38:24]
  always @(posedge clock) begin
    if (reset) begin // @[InstFetch.scala 19:22]
      state <= 2'h0; // @[InstFetch.scala 19:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      state <= 2'h2; // @[InstFetch.scala 45:13]
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (io_stall | io_flush) begin // @[InstFetch.scala 49:19]
        state <= 2'h1;
      end else begin
        state <= 2'h2;
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      state <= _GEN_0;
    end else begin
      state <= _GEN_3;
    end
    if (reset) begin // @[InstFetch.scala 25:19]
      pc <= 32'h30000000; // @[InstFetch.scala 25:19]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(io_stall)) begin // @[InstFetch.scala 48:16]
          pc <= pc_nxt;
        end
      end
    end
    if (reset) begin // @[InstFetch.scala 27:21]
      inst <= 32'h0; // @[InstFetch.scala 27:21]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          inst <= _GEN_4;
        end
      end
    end
    io_out_pc_REG <= ~io_flush; // @[InstFetch.scala 68:50]
    io_out_inst_REG <= ~io_flush; // @[InstFetch.scala 69:52]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  pc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  inst = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_out_pc_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_out_inst_REG = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

module ysyx_210340_Meta(
  input         clock,
  input         reset,
  input  [5:0]  io_idx,
  output [20:0] io_tag_r,
  input  [20:0] io_tag_w,
  input         io_tag_wen,
  output        io_dirty_r,
  input         io_dirty_w,
  input         io_dirty_wen,
  output        io_valid_r,
  input         io_invalidate,
  output        io_dirty_r_async,
  output        io_valid_r_async
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
`endif // RANDOMIZE_REG_INIT
  reg [20:0] tags [0:63]; // @[Cache.scala 38:25]
  wire [20:0] tags_io_tag_r_MPORT_data; // @[Cache.scala 38:25]
  wire [5:0] tags_io_tag_r_MPORT_addr; // @[Cache.scala 38:25]
  wire [20:0] tags_MPORT_data; // @[Cache.scala 38:25]
  wire [5:0] tags_MPORT_addr; // @[Cache.scala 38:25]
  wire  tags_MPORT_mask; // @[Cache.scala 38:25]
  wire  tags_MPORT_en; // @[Cache.scala 38:25]
  reg [5:0] tags_io_tag_r_MPORT_addr_pipe_0;
  reg  valid_0; // @[Cache.scala 40:22]
  reg  valid_1; // @[Cache.scala 40:22]
  reg  valid_2; // @[Cache.scala 40:22]
  reg  valid_3; // @[Cache.scala 40:22]
  reg  valid_4; // @[Cache.scala 40:22]
  reg  valid_5; // @[Cache.scala 40:22]
  reg  valid_6; // @[Cache.scala 40:22]
  reg  valid_7; // @[Cache.scala 40:22]
  reg  valid_8; // @[Cache.scala 40:22]
  reg  valid_9; // @[Cache.scala 40:22]
  reg  valid_10; // @[Cache.scala 40:22]
  reg  valid_11; // @[Cache.scala 40:22]
  reg  valid_12; // @[Cache.scala 40:22]
  reg  valid_13; // @[Cache.scala 40:22]
  reg  valid_14; // @[Cache.scala 40:22]
  reg  valid_15; // @[Cache.scala 40:22]
  reg  valid_16; // @[Cache.scala 40:22]
  reg  valid_17; // @[Cache.scala 40:22]
  reg  valid_18; // @[Cache.scala 40:22]
  reg  valid_19; // @[Cache.scala 40:22]
  reg  valid_20; // @[Cache.scala 40:22]
  reg  valid_21; // @[Cache.scala 40:22]
  reg  valid_22; // @[Cache.scala 40:22]
  reg  valid_23; // @[Cache.scala 40:22]
  reg  valid_24; // @[Cache.scala 40:22]
  reg  valid_25; // @[Cache.scala 40:22]
  reg  valid_26; // @[Cache.scala 40:22]
  reg  valid_27; // @[Cache.scala 40:22]
  reg  valid_28; // @[Cache.scala 40:22]
  reg  valid_29; // @[Cache.scala 40:22]
  reg  valid_30; // @[Cache.scala 40:22]
  reg  valid_31; // @[Cache.scala 40:22]
  reg  valid_32; // @[Cache.scala 40:22]
  reg  valid_33; // @[Cache.scala 40:22]
  reg  valid_34; // @[Cache.scala 40:22]
  reg  valid_35; // @[Cache.scala 40:22]
  reg  valid_36; // @[Cache.scala 40:22]
  reg  valid_37; // @[Cache.scala 40:22]
  reg  valid_38; // @[Cache.scala 40:22]
  reg  valid_39; // @[Cache.scala 40:22]
  reg  valid_40; // @[Cache.scala 40:22]
  reg  valid_41; // @[Cache.scala 40:22]
  reg  valid_42; // @[Cache.scala 40:22]
  reg  valid_43; // @[Cache.scala 40:22]
  reg  valid_44; // @[Cache.scala 40:22]
  reg  valid_45; // @[Cache.scala 40:22]
  reg  valid_46; // @[Cache.scala 40:22]
  reg  valid_47; // @[Cache.scala 40:22]
  reg  valid_48; // @[Cache.scala 40:22]
  reg  valid_49; // @[Cache.scala 40:22]
  reg  valid_50; // @[Cache.scala 40:22]
  reg  valid_51; // @[Cache.scala 40:22]
  reg  valid_52; // @[Cache.scala 40:22]
  reg  valid_53; // @[Cache.scala 40:22]
  reg  valid_54; // @[Cache.scala 40:22]
  reg  valid_55; // @[Cache.scala 40:22]
  reg  valid_56; // @[Cache.scala 40:22]
  reg  valid_57; // @[Cache.scala 40:22]
  reg  valid_58; // @[Cache.scala 40:22]
  reg  valid_59; // @[Cache.scala 40:22]
  reg  valid_60; // @[Cache.scala 40:22]
  reg  valid_61; // @[Cache.scala 40:22]
  reg  valid_62; // @[Cache.scala 40:22]
  reg  valid_63; // @[Cache.scala 40:22]
  reg  dirty_0; // @[Cache.scala 44:22]
  reg  dirty_1; // @[Cache.scala 44:22]
  reg  dirty_2; // @[Cache.scala 44:22]
  reg  dirty_3; // @[Cache.scala 44:22]
  reg  dirty_4; // @[Cache.scala 44:22]
  reg  dirty_5; // @[Cache.scala 44:22]
  reg  dirty_6; // @[Cache.scala 44:22]
  reg  dirty_7; // @[Cache.scala 44:22]
  reg  dirty_8; // @[Cache.scala 44:22]
  reg  dirty_9; // @[Cache.scala 44:22]
  reg  dirty_10; // @[Cache.scala 44:22]
  reg  dirty_11; // @[Cache.scala 44:22]
  reg  dirty_12; // @[Cache.scala 44:22]
  reg  dirty_13; // @[Cache.scala 44:22]
  reg  dirty_14; // @[Cache.scala 44:22]
  reg  dirty_15; // @[Cache.scala 44:22]
  reg  dirty_16; // @[Cache.scala 44:22]
  reg  dirty_17; // @[Cache.scala 44:22]
  reg  dirty_18; // @[Cache.scala 44:22]
  reg  dirty_19; // @[Cache.scala 44:22]
  reg  dirty_20; // @[Cache.scala 44:22]
  reg  dirty_21; // @[Cache.scala 44:22]
  reg  dirty_22; // @[Cache.scala 44:22]
  reg  dirty_23; // @[Cache.scala 44:22]
  reg  dirty_24; // @[Cache.scala 44:22]
  reg  dirty_25; // @[Cache.scala 44:22]
  reg  dirty_26; // @[Cache.scala 44:22]
  reg  dirty_27; // @[Cache.scala 44:22]
  reg  dirty_28; // @[Cache.scala 44:22]
  reg  dirty_29; // @[Cache.scala 44:22]
  reg  dirty_30; // @[Cache.scala 44:22]
  reg  dirty_31; // @[Cache.scala 44:22]
  reg  dirty_32; // @[Cache.scala 44:22]
  reg  dirty_33; // @[Cache.scala 44:22]
  reg  dirty_34; // @[Cache.scala 44:22]
  reg  dirty_35; // @[Cache.scala 44:22]
  reg  dirty_36; // @[Cache.scala 44:22]
  reg  dirty_37; // @[Cache.scala 44:22]
  reg  dirty_38; // @[Cache.scala 44:22]
  reg  dirty_39; // @[Cache.scala 44:22]
  reg  dirty_40; // @[Cache.scala 44:22]
  reg  dirty_41; // @[Cache.scala 44:22]
  reg  dirty_42; // @[Cache.scala 44:22]
  reg  dirty_43; // @[Cache.scala 44:22]
  reg  dirty_44; // @[Cache.scala 44:22]
  reg  dirty_45; // @[Cache.scala 44:22]
  reg  dirty_46; // @[Cache.scala 44:22]
  reg  dirty_47; // @[Cache.scala 44:22]
  reg  dirty_48; // @[Cache.scala 44:22]
  reg  dirty_49; // @[Cache.scala 44:22]
  reg  dirty_50; // @[Cache.scala 44:22]
  reg  dirty_51; // @[Cache.scala 44:22]
  reg  dirty_52; // @[Cache.scala 44:22]
  reg  dirty_53; // @[Cache.scala 44:22]
  reg  dirty_54; // @[Cache.scala 44:22]
  reg  dirty_55; // @[Cache.scala 44:22]
  reg  dirty_56; // @[Cache.scala 44:22]
  reg  dirty_57; // @[Cache.scala 44:22]
  reg  dirty_58; // @[Cache.scala 44:22]
  reg  dirty_59; // @[Cache.scala 44:22]
  reg  dirty_60; // @[Cache.scala 44:22]
  reg  dirty_61; // @[Cache.scala 44:22]
  reg  dirty_62; // @[Cache.scala 44:22]
  reg  dirty_63; // @[Cache.scala 44:22]
  wire  _GEN_0 = 6'h0 == io_idx | valid_0; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_1 = 6'h1 == io_idx | valid_1; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_2 = 6'h2 == io_idx | valid_2; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_3 = 6'h3 == io_idx | valid_3; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_4 = 6'h4 == io_idx | valid_4; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_5 = 6'h5 == io_idx | valid_5; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_6 = 6'h6 == io_idx | valid_6; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_7 = 6'h7 == io_idx | valid_7; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_8 = 6'h8 == io_idx | valid_8; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_9 = 6'h9 == io_idx | valid_9; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_10 = 6'ha == io_idx | valid_10; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_11 = 6'hb == io_idx | valid_11; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_12 = 6'hc == io_idx | valid_12; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_13 = 6'hd == io_idx | valid_13; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_14 = 6'he == io_idx | valid_14; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_15 = 6'hf == io_idx | valid_15; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_16 = 6'h10 == io_idx | valid_16; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_17 = 6'h11 == io_idx | valid_17; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_18 = 6'h12 == io_idx | valid_18; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_19 = 6'h13 == io_idx | valid_19; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_20 = 6'h14 == io_idx | valid_20; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_21 = 6'h15 == io_idx | valid_21; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_22 = 6'h16 == io_idx | valid_22; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_23 = 6'h17 == io_idx | valid_23; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_24 = 6'h18 == io_idx | valid_24; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_25 = 6'h19 == io_idx | valid_25; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_26 = 6'h1a == io_idx | valid_26; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_27 = 6'h1b == io_idx | valid_27; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_28 = 6'h1c == io_idx | valid_28; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_29 = 6'h1d == io_idx | valid_29; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_30 = 6'h1e == io_idx | valid_30; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_31 = 6'h1f == io_idx | valid_31; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_32 = 6'h20 == io_idx | valid_32; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_33 = 6'h21 == io_idx | valid_33; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_34 = 6'h22 == io_idx | valid_34; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_35 = 6'h23 == io_idx | valid_35; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_36 = 6'h24 == io_idx | valid_36; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_37 = 6'h25 == io_idx | valid_37; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_38 = 6'h26 == io_idx | valid_38; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_39 = 6'h27 == io_idx | valid_39; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_40 = 6'h28 == io_idx | valid_40; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_41 = 6'h29 == io_idx | valid_41; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_42 = 6'h2a == io_idx | valid_42; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_43 = 6'h2b == io_idx | valid_43; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_44 = 6'h2c == io_idx | valid_44; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_45 = 6'h2d == io_idx | valid_45; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_46 = 6'h2e == io_idx | valid_46; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_47 = 6'h2f == io_idx | valid_47; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_48 = 6'h30 == io_idx | valid_48; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_49 = 6'h31 == io_idx | valid_49; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_50 = 6'h32 == io_idx | valid_50; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_51 = 6'h33 == io_idx | valid_51; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_52 = 6'h34 == io_idx | valid_52; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_53 = 6'h35 == io_idx | valid_53; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_54 = 6'h36 == io_idx | valid_54; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_55 = 6'h37 == io_idx | valid_55; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_56 = 6'h38 == io_idx | valid_56; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_57 = 6'h39 == io_idx | valid_57; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_58 = 6'h3a == io_idx | valid_58; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_59 = 6'h3b == io_idx | valid_59; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_60 = 6'h3c == io_idx | valid_60; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_61 = 6'h3d == io_idx | valid_61; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_62 = 6'h3e == io_idx | valid_62; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  wire  _GEN_63 = 6'h3f == io_idx | valid_63; // @[Cache.scala 50:16 Cache.scala 50:16 Cache.scala 40:22]
  reg  dirty_r; // @[Cache.scala 55:24]
  wire  _GEN_134 = 6'h1 == io_idx ? dirty_1 : dirty_0; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_135 = 6'h2 == io_idx ? dirty_2 : _GEN_134; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_136 = 6'h3 == io_idx ? dirty_3 : _GEN_135; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_137 = 6'h4 == io_idx ? dirty_4 : _GEN_136; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_138 = 6'h5 == io_idx ? dirty_5 : _GEN_137; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_139 = 6'h6 == io_idx ? dirty_6 : _GEN_138; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_140 = 6'h7 == io_idx ? dirty_7 : _GEN_139; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_141 = 6'h8 == io_idx ? dirty_8 : _GEN_140; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_142 = 6'h9 == io_idx ? dirty_9 : _GEN_141; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_143 = 6'ha == io_idx ? dirty_10 : _GEN_142; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_144 = 6'hb == io_idx ? dirty_11 : _GEN_143; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_145 = 6'hc == io_idx ? dirty_12 : _GEN_144; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_146 = 6'hd == io_idx ? dirty_13 : _GEN_145; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_147 = 6'he == io_idx ? dirty_14 : _GEN_146; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_148 = 6'hf == io_idx ? dirty_15 : _GEN_147; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_149 = 6'h10 == io_idx ? dirty_16 : _GEN_148; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_150 = 6'h11 == io_idx ? dirty_17 : _GEN_149; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_151 = 6'h12 == io_idx ? dirty_18 : _GEN_150; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_152 = 6'h13 == io_idx ? dirty_19 : _GEN_151; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_153 = 6'h14 == io_idx ? dirty_20 : _GEN_152; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_154 = 6'h15 == io_idx ? dirty_21 : _GEN_153; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_155 = 6'h16 == io_idx ? dirty_22 : _GEN_154; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_156 = 6'h17 == io_idx ? dirty_23 : _GEN_155; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_157 = 6'h18 == io_idx ? dirty_24 : _GEN_156; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_158 = 6'h19 == io_idx ? dirty_25 : _GEN_157; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_159 = 6'h1a == io_idx ? dirty_26 : _GEN_158; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_160 = 6'h1b == io_idx ? dirty_27 : _GEN_159; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_161 = 6'h1c == io_idx ? dirty_28 : _GEN_160; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_162 = 6'h1d == io_idx ? dirty_29 : _GEN_161; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_163 = 6'h1e == io_idx ? dirty_30 : _GEN_162; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_164 = 6'h1f == io_idx ? dirty_31 : _GEN_163; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_165 = 6'h20 == io_idx ? dirty_32 : _GEN_164; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_166 = 6'h21 == io_idx ? dirty_33 : _GEN_165; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_167 = 6'h22 == io_idx ? dirty_34 : _GEN_166; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_168 = 6'h23 == io_idx ? dirty_35 : _GEN_167; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_169 = 6'h24 == io_idx ? dirty_36 : _GEN_168; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_170 = 6'h25 == io_idx ? dirty_37 : _GEN_169; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_171 = 6'h26 == io_idx ? dirty_38 : _GEN_170; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_172 = 6'h27 == io_idx ? dirty_39 : _GEN_171; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_173 = 6'h28 == io_idx ? dirty_40 : _GEN_172; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_174 = 6'h29 == io_idx ? dirty_41 : _GEN_173; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_175 = 6'h2a == io_idx ? dirty_42 : _GEN_174; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_176 = 6'h2b == io_idx ? dirty_43 : _GEN_175; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_177 = 6'h2c == io_idx ? dirty_44 : _GEN_176; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_178 = 6'h2d == io_idx ? dirty_45 : _GEN_177; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_179 = 6'h2e == io_idx ? dirty_46 : _GEN_178; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_180 = 6'h2f == io_idx ? dirty_47 : _GEN_179; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_181 = 6'h30 == io_idx ? dirty_48 : _GEN_180; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_182 = 6'h31 == io_idx ? dirty_49 : _GEN_181; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_183 = 6'h32 == io_idx ? dirty_50 : _GEN_182; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_184 = 6'h33 == io_idx ? dirty_51 : _GEN_183; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_185 = 6'h34 == io_idx ? dirty_52 : _GEN_184; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_186 = 6'h35 == io_idx ? dirty_53 : _GEN_185; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_187 = 6'h36 == io_idx ? dirty_54 : _GEN_186; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_188 = 6'h37 == io_idx ? dirty_55 : _GEN_187; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_189 = 6'h38 == io_idx ? dirty_56 : _GEN_188; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_190 = 6'h39 == io_idx ? dirty_57 : _GEN_189; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_191 = 6'h3a == io_idx ? dirty_58 : _GEN_190; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_192 = 6'h3b == io_idx ? dirty_59 : _GEN_191; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_193 = 6'h3c == io_idx ? dirty_60 : _GEN_192; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_194 = 6'h3d == io_idx ? dirty_61 : _GEN_193; // @[Cache.scala 55:24 Cache.scala 55:24]
  wire  _GEN_195 = 6'h3e == io_idx ? dirty_62 : _GEN_194; // @[Cache.scala 55:24 Cache.scala 55:24]
  reg  valid_r; // @[Cache.scala 62:24]
  wire  _GEN_326 = 6'h1 == io_idx ? valid_1 : valid_0; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_327 = 6'h2 == io_idx ? valid_2 : _GEN_326; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_328 = 6'h3 == io_idx ? valid_3 : _GEN_327; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_329 = 6'h4 == io_idx ? valid_4 : _GEN_328; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_330 = 6'h5 == io_idx ? valid_5 : _GEN_329; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_331 = 6'h6 == io_idx ? valid_6 : _GEN_330; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_332 = 6'h7 == io_idx ? valid_7 : _GEN_331; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_333 = 6'h8 == io_idx ? valid_8 : _GEN_332; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_334 = 6'h9 == io_idx ? valid_9 : _GEN_333; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_335 = 6'ha == io_idx ? valid_10 : _GEN_334; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_336 = 6'hb == io_idx ? valid_11 : _GEN_335; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_337 = 6'hc == io_idx ? valid_12 : _GEN_336; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_338 = 6'hd == io_idx ? valid_13 : _GEN_337; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_339 = 6'he == io_idx ? valid_14 : _GEN_338; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_340 = 6'hf == io_idx ? valid_15 : _GEN_339; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_341 = 6'h10 == io_idx ? valid_16 : _GEN_340; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_342 = 6'h11 == io_idx ? valid_17 : _GEN_341; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_343 = 6'h12 == io_idx ? valid_18 : _GEN_342; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_344 = 6'h13 == io_idx ? valid_19 : _GEN_343; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_345 = 6'h14 == io_idx ? valid_20 : _GEN_344; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_346 = 6'h15 == io_idx ? valid_21 : _GEN_345; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_347 = 6'h16 == io_idx ? valid_22 : _GEN_346; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_348 = 6'h17 == io_idx ? valid_23 : _GEN_347; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_349 = 6'h18 == io_idx ? valid_24 : _GEN_348; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_350 = 6'h19 == io_idx ? valid_25 : _GEN_349; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_351 = 6'h1a == io_idx ? valid_26 : _GEN_350; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_352 = 6'h1b == io_idx ? valid_27 : _GEN_351; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_353 = 6'h1c == io_idx ? valid_28 : _GEN_352; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_354 = 6'h1d == io_idx ? valid_29 : _GEN_353; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_355 = 6'h1e == io_idx ? valid_30 : _GEN_354; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_356 = 6'h1f == io_idx ? valid_31 : _GEN_355; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_357 = 6'h20 == io_idx ? valid_32 : _GEN_356; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_358 = 6'h21 == io_idx ? valid_33 : _GEN_357; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_359 = 6'h22 == io_idx ? valid_34 : _GEN_358; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_360 = 6'h23 == io_idx ? valid_35 : _GEN_359; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_361 = 6'h24 == io_idx ? valid_36 : _GEN_360; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_362 = 6'h25 == io_idx ? valid_37 : _GEN_361; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_363 = 6'h26 == io_idx ? valid_38 : _GEN_362; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_364 = 6'h27 == io_idx ? valid_39 : _GEN_363; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_365 = 6'h28 == io_idx ? valid_40 : _GEN_364; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_366 = 6'h29 == io_idx ? valid_41 : _GEN_365; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_367 = 6'h2a == io_idx ? valid_42 : _GEN_366; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_368 = 6'h2b == io_idx ? valid_43 : _GEN_367; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_369 = 6'h2c == io_idx ? valid_44 : _GEN_368; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_370 = 6'h2d == io_idx ? valid_45 : _GEN_369; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_371 = 6'h2e == io_idx ? valid_46 : _GEN_370; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_372 = 6'h2f == io_idx ? valid_47 : _GEN_371; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_373 = 6'h30 == io_idx ? valid_48 : _GEN_372; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_374 = 6'h31 == io_idx ? valid_49 : _GEN_373; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_375 = 6'h32 == io_idx ? valid_50 : _GEN_374; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_376 = 6'h33 == io_idx ? valid_51 : _GEN_375; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_377 = 6'h34 == io_idx ? valid_52 : _GEN_376; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_378 = 6'h35 == io_idx ? valid_53 : _GEN_377; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_379 = 6'h36 == io_idx ? valid_54 : _GEN_378; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_380 = 6'h37 == io_idx ? valid_55 : _GEN_379; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_381 = 6'h38 == io_idx ? valid_56 : _GEN_380; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_382 = 6'h39 == io_idx ? valid_57 : _GEN_381; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_383 = 6'h3a == io_idx ? valid_58 : _GEN_382; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_384 = 6'h3b == io_idx ? valid_59 : _GEN_383; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_385 = 6'h3c == io_idx ? valid_60 : _GEN_384; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_386 = 6'h3d == io_idx ? valid_61 : _GEN_385; // @[Cache.scala 62:24 Cache.scala 62:24]
  wire  _GEN_387 = 6'h3e == io_idx ? valid_62 : _GEN_386; // @[Cache.scala 62:24 Cache.scala 62:24]
  assign tags_io_tag_r_MPORT_addr = tags_io_tag_r_MPORT_addr_pipe_0;
  assign tags_io_tag_r_MPORT_data = tags[tags_io_tag_r_MPORT_addr]; // @[Cache.scala 38:25]
  assign tags_MPORT_data = io_tag_w;
  assign tags_MPORT_addr = io_idx;
  assign tags_MPORT_mask = 1'h1;
  assign tags_MPORT_en = io_tag_wen;
  assign io_tag_r = tags_io_tag_r_MPORT_data; // @[Cache.scala 52:12]
  assign io_dirty_r = dirty_r; // @[Cache.scala 56:14]
  assign io_valid_r = valid_r; // @[Cache.scala 63:14]
  assign io_dirty_r_async = 6'h3f == io_idx ? dirty_63 : _GEN_195; // @[Cache.scala 55:24 Cache.scala 55:24]
  assign io_valid_r_async = 6'h3f == io_idx ? valid_63 : _GEN_387; // @[Cache.scala 62:24 Cache.scala 62:24]
  always @(posedge clock) begin
    if(tags_MPORT_en & tags_MPORT_mask) begin
      tags[tags_MPORT_addr] <= tags_MPORT_data; // @[Cache.scala 38:25]
    end
    tags_io_tag_r_MPORT_addr_pipe_0 <= io_idx;
    if (reset) begin // @[Cache.scala 40:22]
      valid_0 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_0 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_0 <= _GEN_0;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_1 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_1 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_1 <= _GEN_1;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_2 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_2 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_2 <= _GEN_2;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_3 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_3 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_3 <= _GEN_3;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_4 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_4 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_4 <= _GEN_4;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_5 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_5 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_5 <= _GEN_5;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_6 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_6 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_6 <= _GEN_6;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_7 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_7 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_7 <= _GEN_7;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_8 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_8 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_8 <= _GEN_8;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_9 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_9 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_9 <= _GEN_9;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_10 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_10 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_10 <= _GEN_10;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_11 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_11 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_11 <= _GEN_11;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_12 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_12 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_12 <= _GEN_12;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_13 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_13 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_13 <= _GEN_13;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_14 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_14 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_14 <= _GEN_14;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_15 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_15 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_15 <= _GEN_15;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_16 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_16 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_16 <= _GEN_16;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_17 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_17 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_17 <= _GEN_17;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_18 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_18 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_18 <= _GEN_18;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_19 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_19 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_19 <= _GEN_19;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_20 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_20 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_20 <= _GEN_20;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_21 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_21 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_21 <= _GEN_21;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_22 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_22 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_22 <= _GEN_22;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_23 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_23 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_23 <= _GEN_23;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_24 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_24 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_24 <= _GEN_24;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_25 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_25 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_25 <= _GEN_25;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_26 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_26 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_26 <= _GEN_26;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_27 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_27 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_27 <= _GEN_27;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_28 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_28 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_28 <= _GEN_28;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_29 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_29 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_29 <= _GEN_29;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_30 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_30 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_30 <= _GEN_30;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_31 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_31 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_31 <= _GEN_31;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_32 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_32 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_32 <= _GEN_32;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_33 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_33 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_33 <= _GEN_33;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_34 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_34 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_34 <= _GEN_34;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_35 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_35 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_35 <= _GEN_35;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_36 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_36 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_36 <= _GEN_36;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_37 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_37 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_37 <= _GEN_37;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_38 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_38 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_38 <= _GEN_38;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_39 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_39 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_39 <= _GEN_39;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_40 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_40 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_40 <= _GEN_40;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_41 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_41 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_41 <= _GEN_41;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_42 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_42 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_42 <= _GEN_42;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_43 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_43 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_43 <= _GEN_43;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_44 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_44 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_44 <= _GEN_44;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_45 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_45 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_45 <= _GEN_45;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_46 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_46 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_46 <= _GEN_46;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_47 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_47 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_47 <= _GEN_47;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_48 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_48 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_48 <= _GEN_48;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_49 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_49 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_49 <= _GEN_49;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_50 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_50 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_50 <= _GEN_50;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_51 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_51 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_51 <= _GEN_51;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_52 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_52 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_52 <= _GEN_52;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_53 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_53 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_53 <= _GEN_53;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_54 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_54 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_54 <= _GEN_54;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_55 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_55 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_55 <= _GEN_55;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_56 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_56 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_56 <= _GEN_56;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_57 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_57 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_57 <= _GEN_57;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_58 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_58 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_58 <= _GEN_58;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_59 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_59 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_59 <= _GEN_59;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_60 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_60 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_60 <= _GEN_60;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_61 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_61 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_61 <= _GEN_61;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_62 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_62 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_62 <= _GEN_62;
    end
    if (reset) begin // @[Cache.scala 40:22]
      valid_63 <= 1'h0; // @[Cache.scala 40:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      valid_63 <= 1'h0; // @[Cache.scala 68:16]
    end else if (io_tag_wen) begin // @[Cache.scala 48:21]
      valid_63 <= _GEN_63;
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_0 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_0 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h0 == io_idx) begin // @[Cache.scala 59:16]
        dirty_0 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_1 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_1 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h1 == io_idx) begin // @[Cache.scala 59:16]
        dirty_1 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_2 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_2 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h2 == io_idx) begin // @[Cache.scala 59:16]
        dirty_2 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_3 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_3 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h3 == io_idx) begin // @[Cache.scala 59:16]
        dirty_3 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_4 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_4 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h4 == io_idx) begin // @[Cache.scala 59:16]
        dirty_4 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_5 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_5 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h5 == io_idx) begin // @[Cache.scala 59:16]
        dirty_5 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_6 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_6 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h6 == io_idx) begin // @[Cache.scala 59:16]
        dirty_6 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_7 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_7 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h7 == io_idx) begin // @[Cache.scala 59:16]
        dirty_7 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_8 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_8 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h8 == io_idx) begin // @[Cache.scala 59:16]
        dirty_8 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_9 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_9 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h9 == io_idx) begin // @[Cache.scala 59:16]
        dirty_9 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_10 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_10 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'ha == io_idx) begin // @[Cache.scala 59:16]
        dirty_10 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_11 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_11 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'hb == io_idx) begin // @[Cache.scala 59:16]
        dirty_11 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_12 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_12 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'hc == io_idx) begin // @[Cache.scala 59:16]
        dirty_12 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_13 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_13 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'hd == io_idx) begin // @[Cache.scala 59:16]
        dirty_13 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_14 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_14 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'he == io_idx) begin // @[Cache.scala 59:16]
        dirty_14 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_15 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_15 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'hf == io_idx) begin // @[Cache.scala 59:16]
        dirty_15 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_16 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_16 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h10 == io_idx) begin // @[Cache.scala 59:16]
        dirty_16 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_17 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_17 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h11 == io_idx) begin // @[Cache.scala 59:16]
        dirty_17 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_18 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_18 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h12 == io_idx) begin // @[Cache.scala 59:16]
        dirty_18 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_19 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_19 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h13 == io_idx) begin // @[Cache.scala 59:16]
        dirty_19 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_20 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_20 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h14 == io_idx) begin // @[Cache.scala 59:16]
        dirty_20 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_21 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_21 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h15 == io_idx) begin // @[Cache.scala 59:16]
        dirty_21 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_22 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_22 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h16 == io_idx) begin // @[Cache.scala 59:16]
        dirty_22 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_23 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_23 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h17 == io_idx) begin // @[Cache.scala 59:16]
        dirty_23 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_24 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_24 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h18 == io_idx) begin // @[Cache.scala 59:16]
        dirty_24 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_25 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_25 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h19 == io_idx) begin // @[Cache.scala 59:16]
        dirty_25 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_26 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_26 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h1a == io_idx) begin // @[Cache.scala 59:16]
        dirty_26 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_27 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_27 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h1b == io_idx) begin // @[Cache.scala 59:16]
        dirty_27 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_28 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_28 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h1c == io_idx) begin // @[Cache.scala 59:16]
        dirty_28 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_29 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_29 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h1d == io_idx) begin // @[Cache.scala 59:16]
        dirty_29 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_30 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_30 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h1e == io_idx) begin // @[Cache.scala 59:16]
        dirty_30 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_31 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_31 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h1f == io_idx) begin // @[Cache.scala 59:16]
        dirty_31 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_32 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_32 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h20 == io_idx) begin // @[Cache.scala 59:16]
        dirty_32 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_33 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_33 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h21 == io_idx) begin // @[Cache.scala 59:16]
        dirty_33 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_34 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_34 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h22 == io_idx) begin // @[Cache.scala 59:16]
        dirty_34 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_35 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_35 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h23 == io_idx) begin // @[Cache.scala 59:16]
        dirty_35 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_36 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_36 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h24 == io_idx) begin // @[Cache.scala 59:16]
        dirty_36 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_37 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_37 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h25 == io_idx) begin // @[Cache.scala 59:16]
        dirty_37 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_38 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_38 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h26 == io_idx) begin // @[Cache.scala 59:16]
        dirty_38 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_39 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_39 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h27 == io_idx) begin // @[Cache.scala 59:16]
        dirty_39 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_40 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_40 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h28 == io_idx) begin // @[Cache.scala 59:16]
        dirty_40 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_41 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_41 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h29 == io_idx) begin // @[Cache.scala 59:16]
        dirty_41 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_42 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_42 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h2a == io_idx) begin // @[Cache.scala 59:16]
        dirty_42 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_43 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_43 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h2b == io_idx) begin // @[Cache.scala 59:16]
        dirty_43 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_44 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_44 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h2c == io_idx) begin // @[Cache.scala 59:16]
        dirty_44 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_45 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_45 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h2d == io_idx) begin // @[Cache.scala 59:16]
        dirty_45 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_46 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_46 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h2e == io_idx) begin // @[Cache.scala 59:16]
        dirty_46 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_47 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_47 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h2f == io_idx) begin // @[Cache.scala 59:16]
        dirty_47 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_48 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_48 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h30 == io_idx) begin // @[Cache.scala 59:16]
        dirty_48 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_49 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_49 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h31 == io_idx) begin // @[Cache.scala 59:16]
        dirty_49 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_50 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_50 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h32 == io_idx) begin // @[Cache.scala 59:16]
        dirty_50 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_51 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_51 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h33 == io_idx) begin // @[Cache.scala 59:16]
        dirty_51 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_52 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_52 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h34 == io_idx) begin // @[Cache.scala 59:16]
        dirty_52 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_53 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_53 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h35 == io_idx) begin // @[Cache.scala 59:16]
        dirty_53 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_54 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_54 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h36 == io_idx) begin // @[Cache.scala 59:16]
        dirty_54 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_55 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_55 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h37 == io_idx) begin // @[Cache.scala 59:16]
        dirty_55 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_56 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_56 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h38 == io_idx) begin // @[Cache.scala 59:16]
        dirty_56 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_57 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_57 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h39 == io_idx) begin // @[Cache.scala 59:16]
        dirty_57 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_58 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_58 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h3a == io_idx) begin // @[Cache.scala 59:16]
        dirty_58 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_59 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_59 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h3b == io_idx) begin // @[Cache.scala 59:16]
        dirty_59 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_60 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_60 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h3c == io_idx) begin // @[Cache.scala 59:16]
        dirty_60 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_61 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_61 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h3d == io_idx) begin // @[Cache.scala 59:16]
        dirty_61 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_62 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_62 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h3e == io_idx) begin // @[Cache.scala 59:16]
        dirty_62 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (reset) begin // @[Cache.scala 44:22]
      dirty_63 <= 1'h0; // @[Cache.scala 44:22]
    end else if (io_invalidate) begin // @[Cache.scala 65:24]
      dirty_63 <= 1'h0; // @[Cache.scala 67:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 58:23]
      if (6'h3f == io_idx) begin // @[Cache.scala 59:16]
        dirty_63 <= io_dirty_w; // @[Cache.scala 59:16]
      end
    end
    if (6'h3f == io_idx) begin // @[Cache.scala 55:24]
      dirty_r <= dirty_63; // @[Cache.scala 55:24]
    end else if (6'h3e == io_idx) begin // @[Cache.scala 55:24]
      dirty_r <= dirty_62; // @[Cache.scala 55:24]
    end else if (6'h3d == io_idx) begin // @[Cache.scala 55:24]
      dirty_r <= dirty_61; // @[Cache.scala 55:24]
    end else if (6'h3c == io_idx) begin // @[Cache.scala 55:24]
      dirty_r <= dirty_60; // @[Cache.scala 55:24]
    end else begin
      dirty_r <= _GEN_192;
    end
    if (6'h3f == io_idx) begin // @[Cache.scala 62:24]
      valid_r <= valid_63; // @[Cache.scala 62:24]
    end else if (6'h3e == io_idx) begin // @[Cache.scala 62:24]
      valid_r <= valid_62; // @[Cache.scala 62:24]
    end else if (6'h3d == io_idx) begin // @[Cache.scala 62:24]
      valid_r <= valid_61; // @[Cache.scala 62:24]
    end else if (6'h3c == io_idx) begin // @[Cache.scala 62:24]
      valid_r <= valid_60; // @[Cache.scala 62:24]
    end else begin
      valid_r <= _GEN_384;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tags[initvar] = _RAND_0[20:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tags_io_tag_r_MPORT_addr_pipe_0 = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  valid_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  valid_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  valid_3 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  valid_4 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  valid_5 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  valid_6 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  valid_7 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  valid_8 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  valid_9 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  valid_10 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  valid_11 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  valid_12 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  valid_13 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  valid_14 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  valid_15 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  valid_16 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  valid_17 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  valid_18 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  valid_19 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid_20 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  valid_21 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_22 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid_23 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_24 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid_25 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_26 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  valid_27 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  valid_28 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  valid_29 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  valid_30 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  valid_31 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  valid_32 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  valid_33 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  valid_34 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  valid_35 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  valid_36 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  valid_37 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  valid_38 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  valid_39 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  valid_40 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  valid_41 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  valid_42 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  valid_43 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  valid_44 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  valid_45 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  valid_46 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  valid_47 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  valid_48 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  valid_49 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  valid_50 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  valid_51 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  valid_52 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  valid_53 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  valid_54 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  valid_55 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  valid_56 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  valid_57 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  valid_58 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  valid_59 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  valid_60 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  valid_61 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  valid_62 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_63 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  dirty_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  dirty_1 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  dirty_2 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  dirty_3 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  dirty_4 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  dirty_5 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  dirty_6 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  dirty_7 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  dirty_8 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  dirty_9 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  dirty_10 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  dirty_11 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  dirty_12 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  dirty_13 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  dirty_14 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  dirty_15 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  dirty_16 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  dirty_17 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  dirty_18 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  dirty_19 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  dirty_20 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  dirty_21 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  dirty_22 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  dirty_23 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  dirty_24 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  dirty_25 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  dirty_26 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  dirty_27 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  dirty_28 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  dirty_29 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  dirty_30 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  dirty_31 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  dirty_32 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  dirty_33 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  dirty_34 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  dirty_35 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  dirty_36 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  dirty_37 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  dirty_38 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  dirty_39 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  dirty_40 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  dirty_41 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  dirty_42 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  dirty_43 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  dirty_44 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  dirty_45 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  dirty_46 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  dirty_47 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  dirty_48 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  dirty_49 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  dirty_50 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  dirty_51 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  dirty_52 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  dirty_53 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  dirty_54 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  dirty_55 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  dirty_56 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  dirty_57 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  dirty_58 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  dirty_59 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  dirty_60 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  dirty_61 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  dirty_62 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  dirty_63 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  dirty_r = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_r = _RAND_131[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210340_Cache(
  input         clock,
  input         reset,
  output [5:0]   io_sram0_addr,
  output         io_sram0_cen,
  output         io_sram0_wen,
  output [127:0] io_sram0_wdata,
  input  [127:0] io_sram0_rdata,
  output [5:0]   io_sram1_addr,
  output         io_sram1_cen,
  output         io_sram1_wen,
  output [127:0] io_sram1_wdata,
  input  [127:0] io_sram1_rdata,
  output [5:0]   io_sram2_addr,
  output         io_sram2_cen,
  output         io_sram2_wen,
  output [127:0] io_sram2_wdata,
  input  [127:0] io_sram2_rdata,
  output [5:0]   io_sram3_addr,
  output         io_sram3_cen,
  output         io_sram3_wen,
  output [127:0] io_sram3_wdata,
  input  [127:0] io_sram3_rdata,  
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output        io_out_req_bits_aen,
  output        io_out_req_bits_ren,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_req_bits_wlast,
  output        io_out_req_bits_wen,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata,
  input         io_out_resp_bits_rlast,
  input         fence_i_0,
  input         dcache_fi_complete_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [127:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [127:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [63:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [63:0] _RAND_209;
`endif // RANDOMIZE_REG_INIT
  // wire  sram_0_clock; // @[Cache.scala 91:22]
  wire  sram_0_io_en; // @[Cache.scala 91:22]
  wire  sram_0_io_wen; // @[Cache.scala 91:22]
  wire [5:0] sram_0_io_addr; // @[Cache.scala 91:22]
  wire [127:0] sram_0_io_wdata; // @[Cache.scala 91:22]
  wire [127:0] sram_0_io_rdata; // @[Cache.scala 91:22]
  // wire  sram_1_clock; // @[Cache.scala 91:22]
  wire  sram_1_io_en; // @[Cache.scala 91:22]
  wire  sram_1_io_wen; // @[Cache.scala 91:22]
  wire [5:0] sram_1_io_addr; // @[Cache.scala 91:22]
  wire [127:0] sram_1_io_wdata; // @[Cache.scala 91:22]
  wire [127:0] sram_1_io_rdata; // @[Cache.scala 91:22]
  // wire  sram_2_clock; // @[Cache.scala 91:22]
  wire  sram_2_io_en; // @[Cache.scala 91:22]
  wire  sram_2_io_wen; // @[Cache.scala 91:22]
  wire [5:0] sram_2_io_addr; // @[Cache.scala 91:22]
  wire [127:0] sram_2_io_wdata; // @[Cache.scala 91:22]
  wire [127:0] sram_2_io_rdata; // @[Cache.scala 91:22]
  // wire  sram_3_clock; // @[Cache.scala 91:22]
  wire  sram_3_io_en; // @[Cache.scala 91:22]
  wire  sram_3_io_wen; // @[Cache.scala 91:22]
  wire [5:0] sram_3_io_addr; // @[Cache.scala 91:22]
  wire [127:0] sram_3_io_wdata; // @[Cache.scala 91:22]
  wire [127:0] sram_3_io_rdata; // @[Cache.scala 91:22]
  wire  meta_0_clock; // @[Cache.scala 99:22]
  wire  meta_0_reset; // @[Cache.scala 99:22]
  wire [5:0] meta_0_io_idx; // @[Cache.scala 99:22]
  wire [20:0] meta_0_io_tag_r; // @[Cache.scala 99:22]
  wire [20:0] meta_0_io_tag_w; // @[Cache.scala 99:22]
  wire  meta_0_io_tag_wen; // @[Cache.scala 99:22]
  wire  meta_0_io_dirty_r; // @[Cache.scala 99:22]
  wire  meta_0_io_dirty_w; // @[Cache.scala 99:22]
  wire  meta_0_io_dirty_wen; // @[Cache.scala 99:22]
  wire  meta_0_io_valid_r; // @[Cache.scala 99:22]
  wire  meta_0_io_invalidate; // @[Cache.scala 99:22]
  wire  meta_0_io_dirty_r_async; // @[Cache.scala 99:22]
  wire  meta_0_io_valid_r_async; // @[Cache.scala 99:22]
  wire  meta_1_clock; // @[Cache.scala 99:22]
  wire  meta_1_reset; // @[Cache.scala 99:22]
  wire [5:0] meta_1_io_idx; // @[Cache.scala 99:22]
  wire [20:0] meta_1_io_tag_r; // @[Cache.scala 99:22]
  wire [20:0] meta_1_io_tag_w; // @[Cache.scala 99:22]
  wire  meta_1_io_tag_wen; // @[Cache.scala 99:22]
  wire  meta_1_io_dirty_r; // @[Cache.scala 99:22]
  wire  meta_1_io_dirty_w; // @[Cache.scala 99:22]
  wire  meta_1_io_dirty_wen; // @[Cache.scala 99:22]
  wire  meta_1_io_valid_r; // @[Cache.scala 99:22]
  wire  meta_1_io_invalidate; // @[Cache.scala 99:22]
  wire  meta_1_io_dirty_r_async; // @[Cache.scala 99:22]
  wire  meta_1_io_valid_r_async; // @[Cache.scala 99:22]
  wire  meta_2_clock; // @[Cache.scala 99:22]
  wire  meta_2_reset; // @[Cache.scala 99:22]
  wire [5:0] meta_2_io_idx; // @[Cache.scala 99:22]
  wire [20:0] meta_2_io_tag_r; // @[Cache.scala 99:22]
  wire [20:0] meta_2_io_tag_w; // @[Cache.scala 99:22]
  wire  meta_2_io_tag_wen; // @[Cache.scala 99:22]
  wire  meta_2_io_dirty_r; // @[Cache.scala 99:22]
  wire  meta_2_io_dirty_w; // @[Cache.scala 99:22]
  wire  meta_2_io_dirty_wen; // @[Cache.scala 99:22]
  wire  meta_2_io_valid_r; // @[Cache.scala 99:22]
  wire  meta_2_io_invalidate; // @[Cache.scala 99:22]
  wire  meta_2_io_dirty_r_async; // @[Cache.scala 99:22]
  wire  meta_2_io_valid_r_async; // @[Cache.scala 99:22]
  wire  meta_3_clock; // @[Cache.scala 99:22]
  wire  meta_3_reset; // @[Cache.scala 99:22]
  wire [5:0] meta_3_io_idx; // @[Cache.scala 99:22]
  wire [20:0] meta_3_io_tag_r; // @[Cache.scala 99:22]
  wire [20:0] meta_3_io_tag_w; // @[Cache.scala 99:22]
  wire  meta_3_io_tag_wen; // @[Cache.scala 99:22]
  wire  meta_3_io_dirty_r; // @[Cache.scala 99:22]
  wire  meta_3_io_dirty_w; // @[Cache.scala 99:22]
  wire  meta_3_io_dirty_wen; // @[Cache.scala 99:22]
  wire  meta_3_io_valid_r; // @[Cache.scala 99:22]
  wire  meta_3_io_invalidate; // @[Cache.scala 99:22]
  wire  meta_3_io_dirty_r_async; // @[Cache.scala 99:22]
  wire  meta_3_io_valid_r_async; // @[Cache.scala 99:22]
  reg  plru0_0; // @[Cache.scala 131:22]
  reg  plru0_1; // @[Cache.scala 131:22]
  reg  plru0_2; // @[Cache.scala 131:22]
  reg  plru0_3; // @[Cache.scala 131:22]
  reg  plru0_4; // @[Cache.scala 131:22]
  reg  plru0_5; // @[Cache.scala 131:22]
  reg  plru0_6; // @[Cache.scala 131:22]
  reg  plru0_7; // @[Cache.scala 131:22]
  reg  plru0_8; // @[Cache.scala 131:22]
  reg  plru0_9; // @[Cache.scala 131:22]
  reg  plru0_10; // @[Cache.scala 131:22]
  reg  plru0_11; // @[Cache.scala 131:22]
  reg  plru0_12; // @[Cache.scala 131:22]
  reg  plru0_13; // @[Cache.scala 131:22]
  reg  plru0_14; // @[Cache.scala 131:22]
  reg  plru0_15; // @[Cache.scala 131:22]
  reg  plru0_16; // @[Cache.scala 131:22]
  reg  plru0_17; // @[Cache.scala 131:22]
  reg  plru0_18; // @[Cache.scala 131:22]
  reg  plru0_19; // @[Cache.scala 131:22]
  reg  plru0_20; // @[Cache.scala 131:22]
  reg  plru0_21; // @[Cache.scala 131:22]
  reg  plru0_22; // @[Cache.scala 131:22]
  reg  plru0_23; // @[Cache.scala 131:22]
  reg  plru0_24; // @[Cache.scala 131:22]
  reg  plru0_25; // @[Cache.scala 131:22]
  reg  plru0_26; // @[Cache.scala 131:22]
  reg  plru0_27; // @[Cache.scala 131:22]
  reg  plru0_28; // @[Cache.scala 131:22]
  reg  plru0_29; // @[Cache.scala 131:22]
  reg  plru0_30; // @[Cache.scala 131:22]
  reg  plru0_31; // @[Cache.scala 131:22]
  reg  plru0_32; // @[Cache.scala 131:22]
  reg  plru0_33; // @[Cache.scala 131:22]
  reg  plru0_34; // @[Cache.scala 131:22]
  reg  plru0_35; // @[Cache.scala 131:22]
  reg  plru0_36; // @[Cache.scala 131:22]
  reg  plru0_37; // @[Cache.scala 131:22]
  reg  plru0_38; // @[Cache.scala 131:22]
  reg  plru0_39; // @[Cache.scala 131:22]
  reg  plru0_40; // @[Cache.scala 131:22]
  reg  plru0_41; // @[Cache.scala 131:22]
  reg  plru0_42; // @[Cache.scala 131:22]
  reg  plru0_43; // @[Cache.scala 131:22]
  reg  plru0_44; // @[Cache.scala 131:22]
  reg  plru0_45; // @[Cache.scala 131:22]
  reg  plru0_46; // @[Cache.scala 131:22]
  reg  plru0_47; // @[Cache.scala 131:22]
  reg  plru0_48; // @[Cache.scala 131:22]
  reg  plru0_49; // @[Cache.scala 131:22]
  reg  plru0_50; // @[Cache.scala 131:22]
  reg  plru0_51; // @[Cache.scala 131:22]
  reg  plru0_52; // @[Cache.scala 131:22]
  reg  plru0_53; // @[Cache.scala 131:22]
  reg  plru0_54; // @[Cache.scala 131:22]
  reg  plru0_55; // @[Cache.scala 131:22]
  reg  plru0_56; // @[Cache.scala 131:22]
  reg  plru0_57; // @[Cache.scala 131:22]
  reg  plru0_58; // @[Cache.scala 131:22]
  reg  plru0_59; // @[Cache.scala 131:22]
  reg  plru0_60; // @[Cache.scala 131:22]
  reg  plru0_61; // @[Cache.scala 131:22]
  reg  plru0_62; // @[Cache.scala 131:22]
  reg  plru0_63; // @[Cache.scala 131:22]
  reg  plru1_0; // @[Cache.scala 133:22]
  reg  plru1_1; // @[Cache.scala 133:22]
  reg  plru1_2; // @[Cache.scala 133:22]
  reg  plru1_3; // @[Cache.scala 133:22]
  reg  plru1_4; // @[Cache.scala 133:22]
  reg  plru1_5; // @[Cache.scala 133:22]
  reg  plru1_6; // @[Cache.scala 133:22]
  reg  plru1_7; // @[Cache.scala 133:22]
  reg  plru1_8; // @[Cache.scala 133:22]
  reg  plru1_9; // @[Cache.scala 133:22]
  reg  plru1_10; // @[Cache.scala 133:22]
  reg  plru1_11; // @[Cache.scala 133:22]
  reg  plru1_12; // @[Cache.scala 133:22]
  reg  plru1_13; // @[Cache.scala 133:22]
  reg  plru1_14; // @[Cache.scala 133:22]
  reg  plru1_15; // @[Cache.scala 133:22]
  reg  plru1_16; // @[Cache.scala 133:22]
  reg  plru1_17; // @[Cache.scala 133:22]
  reg  plru1_18; // @[Cache.scala 133:22]
  reg  plru1_19; // @[Cache.scala 133:22]
  reg  plru1_20; // @[Cache.scala 133:22]
  reg  plru1_21; // @[Cache.scala 133:22]
  reg  plru1_22; // @[Cache.scala 133:22]
  reg  plru1_23; // @[Cache.scala 133:22]
  reg  plru1_24; // @[Cache.scala 133:22]
  reg  plru1_25; // @[Cache.scala 133:22]
  reg  plru1_26; // @[Cache.scala 133:22]
  reg  plru1_27; // @[Cache.scala 133:22]
  reg  plru1_28; // @[Cache.scala 133:22]
  reg  plru1_29; // @[Cache.scala 133:22]
  reg  plru1_30; // @[Cache.scala 133:22]
  reg  plru1_31; // @[Cache.scala 133:22]
  reg  plru1_32; // @[Cache.scala 133:22]
  reg  plru1_33; // @[Cache.scala 133:22]
  reg  plru1_34; // @[Cache.scala 133:22]
  reg  plru1_35; // @[Cache.scala 133:22]
  reg  plru1_36; // @[Cache.scala 133:22]
  reg  plru1_37; // @[Cache.scala 133:22]
  reg  plru1_38; // @[Cache.scala 133:22]
  reg  plru1_39; // @[Cache.scala 133:22]
  reg  plru1_40; // @[Cache.scala 133:22]
  reg  plru1_41; // @[Cache.scala 133:22]
  reg  plru1_42; // @[Cache.scala 133:22]
  reg  plru1_43; // @[Cache.scala 133:22]
  reg  plru1_44; // @[Cache.scala 133:22]
  reg  plru1_45; // @[Cache.scala 133:22]
  reg  plru1_46; // @[Cache.scala 133:22]
  reg  plru1_47; // @[Cache.scala 133:22]
  reg  plru1_48; // @[Cache.scala 133:22]
  reg  plru1_49; // @[Cache.scala 133:22]
  reg  plru1_50; // @[Cache.scala 133:22]
  reg  plru1_51; // @[Cache.scala 133:22]
  reg  plru1_52; // @[Cache.scala 133:22]
  reg  plru1_53; // @[Cache.scala 133:22]
  reg  plru1_54; // @[Cache.scala 133:22]
  reg  plru1_55; // @[Cache.scala 133:22]
  reg  plru1_56; // @[Cache.scala 133:22]
  reg  plru1_57; // @[Cache.scala 133:22]
  reg  plru1_58; // @[Cache.scala 133:22]
  reg  plru1_59; // @[Cache.scala 133:22]
  reg  plru1_60; // @[Cache.scala 133:22]
  reg  plru1_61; // @[Cache.scala 133:22]
  reg  plru1_62; // @[Cache.scala 133:22]
  reg  plru1_63; // @[Cache.scala 133:22]
  reg  plru2_0; // @[Cache.scala 135:22]
  reg  plru2_1; // @[Cache.scala 135:22]
  reg  plru2_2; // @[Cache.scala 135:22]
  reg  plru2_3; // @[Cache.scala 135:22]
  reg  plru2_4; // @[Cache.scala 135:22]
  reg  plru2_5; // @[Cache.scala 135:22]
  reg  plru2_6; // @[Cache.scala 135:22]
  reg  plru2_7; // @[Cache.scala 135:22]
  reg  plru2_8; // @[Cache.scala 135:22]
  reg  plru2_9; // @[Cache.scala 135:22]
  reg  plru2_10; // @[Cache.scala 135:22]
  reg  plru2_11; // @[Cache.scala 135:22]
  reg  plru2_12; // @[Cache.scala 135:22]
  reg  plru2_13; // @[Cache.scala 135:22]
  reg  plru2_14; // @[Cache.scala 135:22]
  reg  plru2_15; // @[Cache.scala 135:22]
  reg  plru2_16; // @[Cache.scala 135:22]
  reg  plru2_17; // @[Cache.scala 135:22]
  reg  plru2_18; // @[Cache.scala 135:22]
  reg  plru2_19; // @[Cache.scala 135:22]
  reg  plru2_20; // @[Cache.scala 135:22]
  reg  plru2_21; // @[Cache.scala 135:22]
  reg  plru2_22; // @[Cache.scala 135:22]
  reg  plru2_23; // @[Cache.scala 135:22]
  reg  plru2_24; // @[Cache.scala 135:22]
  reg  plru2_25; // @[Cache.scala 135:22]
  reg  plru2_26; // @[Cache.scala 135:22]
  reg  plru2_27; // @[Cache.scala 135:22]
  reg  plru2_28; // @[Cache.scala 135:22]
  reg  plru2_29; // @[Cache.scala 135:22]
  reg  plru2_30; // @[Cache.scala 135:22]
  reg  plru2_31; // @[Cache.scala 135:22]
  reg  plru2_32; // @[Cache.scala 135:22]
  reg  plru2_33; // @[Cache.scala 135:22]
  reg  plru2_34; // @[Cache.scala 135:22]
  reg  plru2_35; // @[Cache.scala 135:22]
  reg  plru2_36; // @[Cache.scala 135:22]
  reg  plru2_37; // @[Cache.scala 135:22]
  reg  plru2_38; // @[Cache.scala 135:22]
  reg  plru2_39; // @[Cache.scala 135:22]
  reg  plru2_40; // @[Cache.scala 135:22]
  reg  plru2_41; // @[Cache.scala 135:22]
  reg  plru2_42; // @[Cache.scala 135:22]
  reg  plru2_43; // @[Cache.scala 135:22]
  reg  plru2_44; // @[Cache.scala 135:22]
  reg  plru2_45; // @[Cache.scala 135:22]
  reg  plru2_46; // @[Cache.scala 135:22]
  reg  plru2_47; // @[Cache.scala 135:22]
  reg  plru2_48; // @[Cache.scala 135:22]
  reg  plru2_49; // @[Cache.scala 135:22]
  reg  plru2_50; // @[Cache.scala 135:22]
  reg  plru2_51; // @[Cache.scala 135:22]
  reg  plru2_52; // @[Cache.scala 135:22]
  reg  plru2_53; // @[Cache.scala 135:22]
  reg  plru2_54; // @[Cache.scala 135:22]
  reg  plru2_55; // @[Cache.scala 135:22]
  reg  plru2_56; // @[Cache.scala 135:22]
  reg  plru2_57; // @[Cache.scala 135:22]
  reg  plru2_58; // @[Cache.scala 135:22]
  reg  plru2_59; // @[Cache.scala 135:22]
  reg  plru2_60; // @[Cache.scala 135:22]
  reg  plru2_61; // @[Cache.scala 135:22]
  reg  plru2_62; // @[Cache.scala 135:22]
  reg  plru2_63; // @[Cache.scala 135:22]
  reg  s2_hit_real_REG; // @[Cache.scala 263:32]
  wire [20:0] tag_out_0 = meta_0_io_tag_r;
  reg [31:0] s2_addr; // @[Cache.scala 209:25]
  wire [20:0] s2_tag = s2_addr[30:10]; // @[Cache.scala 212:25]
  wire  valid_out_0 = meta_0_io_valid_r;
  wire  hit_0 = tag_out_0 == s2_tag & valid_out_0; // @[Cache.scala 222:25]
  wire [20:0] tag_out_1 = meta_1_io_tag_r;
  wire  valid_out_1 = meta_1_io_valid_r;
  wire  hit_1 = tag_out_1 == s2_tag & valid_out_1; // @[Cache.scala 222:25]
  wire [20:0] tag_out_2 = meta_2_io_tag_r;
  wire  valid_out_2 = meta_2_io_valid_r;
  wire  hit_2 = tag_out_2 == s2_tag & valid_out_2; // @[Cache.scala 222:25]
  wire [20:0] tag_out_3 = meta_3_io_tag_r;
  wire  valid_out_3 = meta_3_io_valid_r;
  wire  hit_3 = tag_out_3 == s2_tag & valid_out_3; // @[Cache.scala 222:25]
  wire [3:0] _s2_hit_T = {hit_0,hit_1,hit_2,hit_3}; // @[Cat.scala 30:58]
  wire  s2_hit = |_s2_hit_T; // @[Cache.scala 224:25]
  reg  s2_reg_hit; // @[Cache.scala 231:27]
  wire  s2_hit_real = s2_hit_real_REG ? s2_hit : s2_reg_hit; // @[Cache.scala 263:24]
  reg  s2_wen; // @[Cache.scala 213:25]
  reg [3:0] state; // @[Cache.scala 207:22]
  wire  _hit_ready_T = state == 4'h7; // @[Cache.scala 265:37]
  wire  _hit_ready_T_2 = s2_wen ? state == 4'h7 : state == 4'h0; // @[Cache.scala 265:22]
  wire  hit_ready = s2_hit_real & _hit_ready_T_2; // @[Cache.scala 264:31]
  wire  invalid_ready = state == 4'h8; // @[Cache.scala 267:30]
  wire  fi_ready = (hit_ready | _hit_ready_T) & io_in_resp_ready | invalid_ready; // @[Cache.scala 270:66]
  reg  fi_valid; // @[ID.scala 18:20]
  wire  _GEN_0 = fence_i_0 | fi_valid; // @[ID.scala 24:20 ID.scala 24:24 ID.scala 18:20]
  wire  fi_fire = fi_valid & fi_ready; // @[Cache.scala 163:26]
  wire [5:0] s1_idx = io_in_req_bits_addr[9:4]; // @[Cache.scala 171:25]
  wire [5:0] _GEN_3 = fi_ready ? s1_idx : 6'h0; // @[Cache.scala 181:24 Cache.scala 184:17 Cache.scala 111:15]
  wire  s2_offs = s2_addr[3]; // @[Cache.scala 210:25]
  wire [5:0] s2_idx = s2_addr[9:4]; // @[Cache.scala 211:25]
  reg [63:0] s2_wdata; // @[Cache.scala 214:25]
  reg [7:0] s2_wmask; // @[Cache.scala 215:25]
  wire [3:0] _s2_way_T = {hit_3,hit_2,hit_1,hit_0}; // @[OneHot.scala 22:45]
  wire [1:0] s2_way_hi_1 = _s2_way_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] s2_way_lo_1 = _s2_way_T[1:0]; // @[OneHot.scala 31:18]
  wire  s2_way_hi_2 = |s2_way_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _s2_way_T_1 = s2_way_hi_1 | s2_way_lo_1; // @[OneHot.scala 32:28]
  wire  s2_way_lo_2 = _s2_way_T_1[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] s2_way = {s2_way_hi_2,s2_way_lo_2}; // @[Cat.scala 30:58]
  reg [127:0] s2_reg_rdata; // @[Cache.scala 233:29]
  reg  s2_reg_dirty; // @[Cache.scala 234:29]
  reg [20:0] s2_reg_tag_r; // @[Cache.scala 235:29]
  reg [127:0] s2_reg_dat_w; // @[Cache.scala 236:29]
  reg  REG; // @[Cache.scala 244:41]
  wire [127:0] sram_out_0 = sram_0_io_rdata;
  wire [127:0] sram_out_1 = sram_1_io_rdata;
  wire [127:0] _GEN_5 = 2'h1 == s2_way ? sram_out_1 : sram_out_0; // @[Cache.scala 249:18 Cache.scala 249:18]
  wire [127:0] sram_out_2 = sram_2_io_rdata;
  wire [127:0] _GEN_6 = 2'h2 == s2_way ? sram_out_2 : _GEN_5; // @[Cache.scala 249:18 Cache.scala 249:18]
  wire [127:0] sram_out_3 = sram_3_io_rdata;
  wire [127:0] _GEN_7 = 2'h3 == s2_way ? sram_out_3 : _GEN_6; // @[Cache.scala 249:18 Cache.scala 249:18]
  wire  _GEN_37 = 6'h1 == s2_idx ? plru0_1 : plru0_0; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_38 = 6'h2 == s2_idx ? plru0_2 : _GEN_37; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_39 = 6'h3 == s2_idx ? plru0_3 : _GEN_38; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_40 = 6'h4 == s2_idx ? plru0_4 : _GEN_39; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_41 = 6'h5 == s2_idx ? plru0_5 : _GEN_40; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_42 = 6'h6 == s2_idx ? plru0_6 : _GEN_41; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_43 = 6'h7 == s2_idx ? plru0_7 : _GEN_42; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_44 = 6'h8 == s2_idx ? plru0_8 : _GEN_43; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_45 = 6'h9 == s2_idx ? plru0_9 : _GEN_44; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_46 = 6'ha == s2_idx ? plru0_10 : _GEN_45; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_47 = 6'hb == s2_idx ? plru0_11 : _GEN_46; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_48 = 6'hc == s2_idx ? plru0_12 : _GEN_47; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_49 = 6'hd == s2_idx ? plru0_13 : _GEN_48; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_50 = 6'he == s2_idx ? plru0_14 : _GEN_49; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_51 = 6'hf == s2_idx ? plru0_15 : _GEN_50; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_52 = 6'h10 == s2_idx ? plru0_16 : _GEN_51; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_53 = 6'h11 == s2_idx ? plru0_17 : _GEN_52; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_54 = 6'h12 == s2_idx ? plru0_18 : _GEN_53; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_55 = 6'h13 == s2_idx ? plru0_19 : _GEN_54; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_56 = 6'h14 == s2_idx ? plru0_20 : _GEN_55; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_57 = 6'h15 == s2_idx ? plru0_21 : _GEN_56; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_58 = 6'h16 == s2_idx ? plru0_22 : _GEN_57; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_59 = 6'h17 == s2_idx ? plru0_23 : _GEN_58; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_60 = 6'h18 == s2_idx ? plru0_24 : _GEN_59; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_61 = 6'h19 == s2_idx ? plru0_25 : _GEN_60; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_62 = 6'h1a == s2_idx ? plru0_26 : _GEN_61; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_63 = 6'h1b == s2_idx ? plru0_27 : _GEN_62; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_64 = 6'h1c == s2_idx ? plru0_28 : _GEN_63; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_65 = 6'h1d == s2_idx ? plru0_29 : _GEN_64; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_66 = 6'h1e == s2_idx ? plru0_30 : _GEN_65; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_67 = 6'h1f == s2_idx ? plru0_31 : _GEN_66; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_68 = 6'h20 == s2_idx ? plru0_32 : _GEN_67; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_69 = 6'h21 == s2_idx ? plru0_33 : _GEN_68; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_70 = 6'h22 == s2_idx ? plru0_34 : _GEN_69; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_71 = 6'h23 == s2_idx ? plru0_35 : _GEN_70; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_72 = 6'h24 == s2_idx ? plru0_36 : _GEN_71; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_73 = 6'h25 == s2_idx ? plru0_37 : _GEN_72; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_74 = 6'h26 == s2_idx ? plru0_38 : _GEN_73; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_75 = 6'h27 == s2_idx ? plru0_39 : _GEN_74; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_76 = 6'h28 == s2_idx ? plru0_40 : _GEN_75; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_77 = 6'h29 == s2_idx ? plru0_41 : _GEN_76; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_78 = 6'h2a == s2_idx ? plru0_42 : _GEN_77; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_79 = 6'h2b == s2_idx ? plru0_43 : _GEN_78; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_80 = 6'h2c == s2_idx ? plru0_44 : _GEN_79; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_81 = 6'h2d == s2_idx ? plru0_45 : _GEN_80; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_82 = 6'h2e == s2_idx ? plru0_46 : _GEN_81; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_83 = 6'h2f == s2_idx ? plru0_47 : _GEN_82; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_84 = 6'h30 == s2_idx ? plru0_48 : _GEN_83; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_85 = 6'h31 == s2_idx ? plru0_49 : _GEN_84; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_86 = 6'h32 == s2_idx ? plru0_50 : _GEN_85; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_87 = 6'h33 == s2_idx ? plru0_51 : _GEN_86; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_88 = 6'h34 == s2_idx ? plru0_52 : _GEN_87; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_89 = 6'h35 == s2_idx ? plru0_53 : _GEN_88; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_90 = 6'h36 == s2_idx ? plru0_54 : _GEN_89; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_91 = 6'h37 == s2_idx ? plru0_55 : _GEN_90; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_92 = 6'h38 == s2_idx ? plru0_56 : _GEN_91; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_93 = 6'h39 == s2_idx ? plru0_57 : _GEN_92; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_94 = 6'h3a == s2_idx ? plru0_58 : _GEN_93; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_95 = 6'h3b == s2_idx ? plru0_59 : _GEN_94; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_96 = 6'h3c == s2_idx ? plru0_60 : _GEN_95; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_97 = 6'h3d == s2_idx ? plru0_61 : _GEN_96; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_98 = 6'h3e == s2_idx ? plru0_62 : _GEN_97; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_99 = 6'h3f == s2_idx ? plru0_63 : _GEN_98; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_101 = 6'h1 == s2_idx ? plru1_1 : plru1_0; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_102 = 6'h2 == s2_idx ? plru1_2 : _GEN_101; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_103 = 6'h3 == s2_idx ? plru1_3 : _GEN_102; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_104 = 6'h4 == s2_idx ? plru1_4 : _GEN_103; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_105 = 6'h5 == s2_idx ? plru1_5 : _GEN_104; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_106 = 6'h6 == s2_idx ? plru1_6 : _GEN_105; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_107 = 6'h7 == s2_idx ? plru1_7 : _GEN_106; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_108 = 6'h8 == s2_idx ? plru1_8 : _GEN_107; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_109 = 6'h9 == s2_idx ? plru1_9 : _GEN_108; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_110 = 6'ha == s2_idx ? plru1_10 : _GEN_109; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_111 = 6'hb == s2_idx ? plru1_11 : _GEN_110; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_112 = 6'hc == s2_idx ? plru1_12 : _GEN_111; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_113 = 6'hd == s2_idx ? plru1_13 : _GEN_112; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_114 = 6'he == s2_idx ? plru1_14 : _GEN_113; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_115 = 6'hf == s2_idx ? plru1_15 : _GEN_114; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_116 = 6'h10 == s2_idx ? plru1_16 : _GEN_115; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_117 = 6'h11 == s2_idx ? plru1_17 : _GEN_116; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_118 = 6'h12 == s2_idx ? plru1_18 : _GEN_117; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_119 = 6'h13 == s2_idx ? plru1_19 : _GEN_118; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_120 = 6'h14 == s2_idx ? plru1_20 : _GEN_119; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_121 = 6'h15 == s2_idx ? plru1_21 : _GEN_120; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_122 = 6'h16 == s2_idx ? plru1_22 : _GEN_121; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_123 = 6'h17 == s2_idx ? plru1_23 : _GEN_122; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_124 = 6'h18 == s2_idx ? plru1_24 : _GEN_123; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_125 = 6'h19 == s2_idx ? plru1_25 : _GEN_124; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_126 = 6'h1a == s2_idx ? plru1_26 : _GEN_125; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_127 = 6'h1b == s2_idx ? plru1_27 : _GEN_126; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_128 = 6'h1c == s2_idx ? plru1_28 : _GEN_127; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_129 = 6'h1d == s2_idx ? plru1_29 : _GEN_128; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_130 = 6'h1e == s2_idx ? plru1_30 : _GEN_129; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_131 = 6'h1f == s2_idx ? plru1_31 : _GEN_130; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_132 = 6'h20 == s2_idx ? plru1_32 : _GEN_131; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_133 = 6'h21 == s2_idx ? plru1_33 : _GEN_132; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_134 = 6'h22 == s2_idx ? plru1_34 : _GEN_133; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_135 = 6'h23 == s2_idx ? plru1_35 : _GEN_134; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_136 = 6'h24 == s2_idx ? plru1_36 : _GEN_135; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_137 = 6'h25 == s2_idx ? plru1_37 : _GEN_136; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_138 = 6'h26 == s2_idx ? plru1_38 : _GEN_137; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_139 = 6'h27 == s2_idx ? plru1_39 : _GEN_138; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_140 = 6'h28 == s2_idx ? plru1_40 : _GEN_139; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_141 = 6'h29 == s2_idx ? plru1_41 : _GEN_140; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_142 = 6'h2a == s2_idx ? plru1_42 : _GEN_141; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_143 = 6'h2b == s2_idx ? plru1_43 : _GEN_142; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_144 = 6'h2c == s2_idx ? plru1_44 : _GEN_143; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_145 = 6'h2d == s2_idx ? plru1_45 : _GEN_144; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_146 = 6'h2e == s2_idx ? plru1_46 : _GEN_145; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_147 = 6'h2f == s2_idx ? plru1_47 : _GEN_146; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_148 = 6'h30 == s2_idx ? plru1_48 : _GEN_147; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_149 = 6'h31 == s2_idx ? plru1_49 : _GEN_148; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_150 = 6'h32 == s2_idx ? plru1_50 : _GEN_149; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_151 = 6'h33 == s2_idx ? plru1_51 : _GEN_150; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_152 = 6'h34 == s2_idx ? plru1_52 : _GEN_151; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_153 = 6'h35 == s2_idx ? plru1_53 : _GEN_152; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_154 = 6'h36 == s2_idx ? plru1_54 : _GEN_153; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_155 = 6'h37 == s2_idx ? plru1_55 : _GEN_154; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_156 = 6'h38 == s2_idx ? plru1_56 : _GEN_155; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_157 = 6'h39 == s2_idx ? plru1_57 : _GEN_156; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_158 = 6'h3a == s2_idx ? plru1_58 : _GEN_157; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_159 = 6'h3b == s2_idx ? plru1_59 : _GEN_158; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_160 = 6'h3c == s2_idx ? plru1_60 : _GEN_159; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_161 = 6'h3d == s2_idx ? plru1_61 : _GEN_160; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_162 = 6'h3e == s2_idx ? plru1_62 : _GEN_161; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_163 = 6'h3f == s2_idx ? plru1_63 : _GEN_162; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_165 = 6'h1 == s2_idx ? plru2_1 : plru2_0; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_166 = 6'h2 == s2_idx ? plru2_2 : _GEN_165; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_167 = 6'h3 == s2_idx ? plru2_3 : _GEN_166; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_168 = 6'h4 == s2_idx ? plru2_4 : _GEN_167; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_169 = 6'h5 == s2_idx ? plru2_5 : _GEN_168; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_170 = 6'h6 == s2_idx ? plru2_6 : _GEN_169; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_171 = 6'h7 == s2_idx ? plru2_7 : _GEN_170; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_172 = 6'h8 == s2_idx ? plru2_8 : _GEN_171; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_173 = 6'h9 == s2_idx ? plru2_9 : _GEN_172; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_174 = 6'ha == s2_idx ? plru2_10 : _GEN_173; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_175 = 6'hb == s2_idx ? plru2_11 : _GEN_174; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_176 = 6'hc == s2_idx ? plru2_12 : _GEN_175; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_177 = 6'hd == s2_idx ? plru2_13 : _GEN_176; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_178 = 6'he == s2_idx ? plru2_14 : _GEN_177; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_179 = 6'hf == s2_idx ? plru2_15 : _GEN_178; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_180 = 6'h10 == s2_idx ? plru2_16 : _GEN_179; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_181 = 6'h11 == s2_idx ? plru2_17 : _GEN_180; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_182 = 6'h12 == s2_idx ? plru2_18 : _GEN_181; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_183 = 6'h13 == s2_idx ? plru2_19 : _GEN_182; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_184 = 6'h14 == s2_idx ? plru2_20 : _GEN_183; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_185 = 6'h15 == s2_idx ? plru2_21 : _GEN_184; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_186 = 6'h16 == s2_idx ? plru2_22 : _GEN_185; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_187 = 6'h17 == s2_idx ? plru2_23 : _GEN_186; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_188 = 6'h18 == s2_idx ? plru2_24 : _GEN_187; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_189 = 6'h19 == s2_idx ? plru2_25 : _GEN_188; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_190 = 6'h1a == s2_idx ? plru2_26 : _GEN_189; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_191 = 6'h1b == s2_idx ? plru2_27 : _GEN_190; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_192 = 6'h1c == s2_idx ? plru2_28 : _GEN_191; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_193 = 6'h1d == s2_idx ? plru2_29 : _GEN_192; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_194 = 6'h1e == s2_idx ? plru2_30 : _GEN_193; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_195 = 6'h1f == s2_idx ? plru2_31 : _GEN_194; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_196 = 6'h20 == s2_idx ? plru2_32 : _GEN_195; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_197 = 6'h21 == s2_idx ? plru2_33 : _GEN_196; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_198 = 6'h22 == s2_idx ? plru2_34 : _GEN_197; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_199 = 6'h23 == s2_idx ? plru2_35 : _GEN_198; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_200 = 6'h24 == s2_idx ? plru2_36 : _GEN_199; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_201 = 6'h25 == s2_idx ? plru2_37 : _GEN_200; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_202 = 6'h26 == s2_idx ? plru2_38 : _GEN_201; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_203 = 6'h27 == s2_idx ? plru2_39 : _GEN_202; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_204 = 6'h28 == s2_idx ? plru2_40 : _GEN_203; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_205 = 6'h29 == s2_idx ? plru2_41 : _GEN_204; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_206 = 6'h2a == s2_idx ? plru2_42 : _GEN_205; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_207 = 6'h2b == s2_idx ? plru2_43 : _GEN_206; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_208 = 6'h2c == s2_idx ? plru2_44 : _GEN_207; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_209 = 6'h2d == s2_idx ? plru2_45 : _GEN_208; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_210 = 6'h2e == s2_idx ? plru2_46 : _GEN_209; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_211 = 6'h2f == s2_idx ? plru2_47 : _GEN_210; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_212 = 6'h30 == s2_idx ? plru2_48 : _GEN_211; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_213 = 6'h31 == s2_idx ? plru2_49 : _GEN_212; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_214 = 6'h32 == s2_idx ? plru2_50 : _GEN_213; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_215 = 6'h33 == s2_idx ? plru2_51 : _GEN_214; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_216 = 6'h34 == s2_idx ? plru2_52 : _GEN_215; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_217 = 6'h35 == s2_idx ? plru2_53 : _GEN_216; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_218 = 6'h36 == s2_idx ? plru2_54 : _GEN_217; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_219 = 6'h37 == s2_idx ? plru2_55 : _GEN_218; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_220 = 6'h38 == s2_idx ? plru2_56 : _GEN_219; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_221 = 6'h39 == s2_idx ? plru2_57 : _GEN_220; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_222 = 6'h3a == s2_idx ? plru2_58 : _GEN_221; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_223 = 6'h3b == s2_idx ? plru2_59 : _GEN_222; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_224 = 6'h3c == s2_idx ? plru2_60 : _GEN_223; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_225 = 6'h3d == s2_idx ? plru2_61 : _GEN_224; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_226 = 6'h3e == s2_idx ? plru2_62 : _GEN_225; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_227 = 6'h3f == s2_idx ? plru2_63 : _GEN_226; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  replace_way_lo = ~_GEN_99 ? _GEN_163 : _GEN_227; // @[Cache.scala 256:25]
  wire [1:0] replace_way = {_GEN_99,replace_way_lo}; // @[Cat.scala 30:58]
  wire  dirty_out_0 = meta_0_io_dirty_r;
  wire  dirty_out_1 = meta_1_io_dirty_r;
  wire  _GEN_9 = 2'h1 == replace_way ? dirty_out_1 : dirty_out_0; // @[Cache.scala 250:18 Cache.scala 250:18]
  wire  dirty_out_2 = meta_2_io_dirty_r;
  wire  _GEN_10 = 2'h2 == replace_way ? dirty_out_2 : _GEN_9; // @[Cache.scala 250:18 Cache.scala 250:18]
  wire  dirty_out_3 = meta_3_io_dirty_r;
  wire [20:0] _GEN_13 = 2'h1 == replace_way ? tag_out_1 : tag_out_0; // @[Cache.scala 251:18 Cache.scala 251:18]
  wire [20:0] _GEN_14 = 2'h2 == replace_way ? tag_out_2 : _GEN_13; // @[Cache.scala 251:18 Cache.scala 251:18]
  wire [127:0] _GEN_17 = 2'h1 == replace_way ? sram_out_1 : sram_out_0; // @[Cache.scala 252:18 Cache.scala 252:18]
  wire [127:0] _GEN_18 = 2'h2 == replace_way ? sram_out_2 : _GEN_17; // @[Cache.scala 252:18 Cache.scala 252:18]
  wire  _GEN_27 = fi_ready ? io_in_req_bits_wen : s2_wen; // @[Cache.scala 238:24 Cache.scala 241:14 Cache.scala 213:25]
  reg [63:0] wdata1; // @[Cache.scala 258:23]
  reg [63:0] wdata2; // @[Cache.scala 259:23]
  wire  _T_2 = 4'h0 == state; // @[Conditional.scala 37:30]
  reg  REG_1; // @[Cache.scala 284:20]
  wire [63:0] _io_in_resp_bits_rdata_T_3 = s2_offs ? _GEN_7[127:64] : _GEN_7[63:0]; // @[Cache.scala 285:34]
  wire [63:0] _io_in_resp_bits_rdata_T_7 = s2_offs ? s2_reg_rdata[127:64] : s2_reg_rdata[63:0]; // @[Cache.scala 287:34]
  wire [63:0] _GEN_228 = REG_1 ? _io_in_resp_bits_rdata_T_3 : _io_in_resp_bits_rdata_T_7; // @[Cache.scala 284:37 Cache.scala 285:28 Cache.scala 287:28]
  reg  REG_2; // @[Cache.scala 289:20]
  wire  _plru0_T_1 = ~s2_way[1]; // @[Cache.scala 138:19]
  wire  _GEN_229 = 6'h0 == s2_idx ? ~s2_way[1] : plru0_0; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_230 = 6'h1 == s2_idx ? ~s2_way[1] : plru0_1; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_231 = 6'h2 == s2_idx ? ~s2_way[1] : plru0_2; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_232 = 6'h3 == s2_idx ? ~s2_way[1] : plru0_3; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_233 = 6'h4 == s2_idx ? ~s2_way[1] : plru0_4; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_234 = 6'h5 == s2_idx ? ~s2_way[1] : plru0_5; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_235 = 6'h6 == s2_idx ? ~s2_way[1] : plru0_6; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_236 = 6'h7 == s2_idx ? ~s2_way[1] : plru0_7; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_237 = 6'h8 == s2_idx ? ~s2_way[1] : plru0_8; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_238 = 6'h9 == s2_idx ? ~s2_way[1] : plru0_9; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_239 = 6'ha == s2_idx ? ~s2_way[1] : plru0_10; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_240 = 6'hb == s2_idx ? ~s2_way[1] : plru0_11; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_241 = 6'hc == s2_idx ? ~s2_way[1] : plru0_12; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_242 = 6'hd == s2_idx ? ~s2_way[1] : plru0_13; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_243 = 6'he == s2_idx ? ~s2_way[1] : plru0_14; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_244 = 6'hf == s2_idx ? ~s2_way[1] : plru0_15; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_245 = 6'h10 == s2_idx ? ~s2_way[1] : plru0_16; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_246 = 6'h11 == s2_idx ? ~s2_way[1] : plru0_17; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_247 = 6'h12 == s2_idx ? ~s2_way[1] : plru0_18; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_248 = 6'h13 == s2_idx ? ~s2_way[1] : plru0_19; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_249 = 6'h14 == s2_idx ? ~s2_way[1] : plru0_20; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_250 = 6'h15 == s2_idx ? ~s2_way[1] : plru0_21; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_251 = 6'h16 == s2_idx ? ~s2_way[1] : plru0_22; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_252 = 6'h17 == s2_idx ? ~s2_way[1] : plru0_23; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_253 = 6'h18 == s2_idx ? ~s2_way[1] : plru0_24; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_254 = 6'h19 == s2_idx ? ~s2_way[1] : plru0_25; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_255 = 6'h1a == s2_idx ? ~s2_way[1] : plru0_26; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_256 = 6'h1b == s2_idx ? ~s2_way[1] : plru0_27; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_257 = 6'h1c == s2_idx ? ~s2_way[1] : plru0_28; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_258 = 6'h1d == s2_idx ? ~s2_way[1] : plru0_29; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_259 = 6'h1e == s2_idx ? ~s2_way[1] : plru0_30; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_260 = 6'h1f == s2_idx ? ~s2_way[1] : plru0_31; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_261 = 6'h20 == s2_idx ? ~s2_way[1] : plru0_32; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_262 = 6'h21 == s2_idx ? ~s2_way[1] : plru0_33; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_263 = 6'h22 == s2_idx ? ~s2_way[1] : plru0_34; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_264 = 6'h23 == s2_idx ? ~s2_way[1] : plru0_35; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_265 = 6'h24 == s2_idx ? ~s2_way[1] : plru0_36; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_266 = 6'h25 == s2_idx ? ~s2_way[1] : plru0_37; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_267 = 6'h26 == s2_idx ? ~s2_way[1] : plru0_38; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_268 = 6'h27 == s2_idx ? ~s2_way[1] : plru0_39; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_269 = 6'h28 == s2_idx ? ~s2_way[1] : plru0_40; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_270 = 6'h29 == s2_idx ? ~s2_way[1] : plru0_41; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_271 = 6'h2a == s2_idx ? ~s2_way[1] : plru0_42; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_272 = 6'h2b == s2_idx ? ~s2_way[1] : plru0_43; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_273 = 6'h2c == s2_idx ? ~s2_way[1] : plru0_44; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_274 = 6'h2d == s2_idx ? ~s2_way[1] : plru0_45; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_275 = 6'h2e == s2_idx ? ~s2_way[1] : plru0_46; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_276 = 6'h2f == s2_idx ? ~s2_way[1] : plru0_47; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_277 = 6'h30 == s2_idx ? ~s2_way[1] : plru0_48; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_278 = 6'h31 == s2_idx ? ~s2_way[1] : plru0_49; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_279 = 6'h32 == s2_idx ? ~s2_way[1] : plru0_50; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_280 = 6'h33 == s2_idx ? ~s2_way[1] : plru0_51; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_281 = 6'h34 == s2_idx ? ~s2_way[1] : plru0_52; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_282 = 6'h35 == s2_idx ? ~s2_way[1] : plru0_53; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_283 = 6'h36 == s2_idx ? ~s2_way[1] : plru0_54; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_284 = 6'h37 == s2_idx ? ~s2_way[1] : plru0_55; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_285 = 6'h38 == s2_idx ? ~s2_way[1] : plru0_56; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_286 = 6'h39 == s2_idx ? ~s2_way[1] : plru0_57; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_287 = 6'h3a == s2_idx ? ~s2_way[1] : plru0_58; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_288 = 6'h3b == s2_idx ? ~s2_way[1] : plru0_59; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_289 = 6'h3c == s2_idx ? ~s2_way[1] : plru0_60; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_290 = 6'h3d == s2_idx ? ~s2_way[1] : plru0_61; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_291 = 6'h3e == s2_idx ? ~s2_way[1] : plru0_62; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_292 = 6'h3f == s2_idx ? ~s2_way[1] : plru0_63; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _plru1_T_1 = ~s2_way[0]; // @[Cache.scala 140:21]
  wire  _GEN_293 = 6'h0 == s2_idx ? ~s2_way[0] : plru1_0; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_294 = 6'h1 == s2_idx ? ~s2_way[0] : plru1_1; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_295 = 6'h2 == s2_idx ? ~s2_way[0] : plru1_2; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_296 = 6'h3 == s2_idx ? ~s2_way[0] : plru1_3; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_297 = 6'h4 == s2_idx ? ~s2_way[0] : plru1_4; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_298 = 6'h5 == s2_idx ? ~s2_way[0] : plru1_5; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_299 = 6'h6 == s2_idx ? ~s2_way[0] : plru1_6; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_300 = 6'h7 == s2_idx ? ~s2_way[0] : plru1_7; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_301 = 6'h8 == s2_idx ? ~s2_way[0] : plru1_8; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_302 = 6'h9 == s2_idx ? ~s2_way[0] : plru1_9; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_303 = 6'ha == s2_idx ? ~s2_way[0] : plru1_10; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_304 = 6'hb == s2_idx ? ~s2_way[0] : plru1_11; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_305 = 6'hc == s2_idx ? ~s2_way[0] : plru1_12; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_306 = 6'hd == s2_idx ? ~s2_way[0] : plru1_13; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_307 = 6'he == s2_idx ? ~s2_way[0] : plru1_14; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_308 = 6'hf == s2_idx ? ~s2_way[0] : plru1_15; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_309 = 6'h10 == s2_idx ? ~s2_way[0] : plru1_16; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_310 = 6'h11 == s2_idx ? ~s2_way[0] : plru1_17; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_311 = 6'h12 == s2_idx ? ~s2_way[0] : plru1_18; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_312 = 6'h13 == s2_idx ? ~s2_way[0] : plru1_19; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_313 = 6'h14 == s2_idx ? ~s2_way[0] : plru1_20; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_314 = 6'h15 == s2_idx ? ~s2_way[0] : plru1_21; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_315 = 6'h16 == s2_idx ? ~s2_way[0] : plru1_22; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_316 = 6'h17 == s2_idx ? ~s2_way[0] : plru1_23; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_317 = 6'h18 == s2_idx ? ~s2_way[0] : plru1_24; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_318 = 6'h19 == s2_idx ? ~s2_way[0] : plru1_25; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_319 = 6'h1a == s2_idx ? ~s2_way[0] : plru1_26; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_320 = 6'h1b == s2_idx ? ~s2_way[0] : plru1_27; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_321 = 6'h1c == s2_idx ? ~s2_way[0] : plru1_28; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_322 = 6'h1d == s2_idx ? ~s2_way[0] : plru1_29; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_323 = 6'h1e == s2_idx ? ~s2_way[0] : plru1_30; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_324 = 6'h1f == s2_idx ? ~s2_way[0] : plru1_31; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_325 = 6'h20 == s2_idx ? ~s2_way[0] : plru1_32; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_326 = 6'h21 == s2_idx ? ~s2_way[0] : plru1_33; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_327 = 6'h22 == s2_idx ? ~s2_way[0] : plru1_34; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_328 = 6'h23 == s2_idx ? ~s2_way[0] : plru1_35; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_329 = 6'h24 == s2_idx ? ~s2_way[0] : plru1_36; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_330 = 6'h25 == s2_idx ? ~s2_way[0] : plru1_37; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_331 = 6'h26 == s2_idx ? ~s2_way[0] : plru1_38; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_332 = 6'h27 == s2_idx ? ~s2_way[0] : plru1_39; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_333 = 6'h28 == s2_idx ? ~s2_way[0] : plru1_40; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_334 = 6'h29 == s2_idx ? ~s2_way[0] : plru1_41; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_335 = 6'h2a == s2_idx ? ~s2_way[0] : plru1_42; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_336 = 6'h2b == s2_idx ? ~s2_way[0] : plru1_43; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_337 = 6'h2c == s2_idx ? ~s2_way[0] : plru1_44; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_338 = 6'h2d == s2_idx ? ~s2_way[0] : plru1_45; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_339 = 6'h2e == s2_idx ? ~s2_way[0] : plru1_46; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_340 = 6'h2f == s2_idx ? ~s2_way[0] : plru1_47; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_341 = 6'h30 == s2_idx ? ~s2_way[0] : plru1_48; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_342 = 6'h31 == s2_idx ? ~s2_way[0] : plru1_49; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_343 = 6'h32 == s2_idx ? ~s2_way[0] : plru1_50; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_344 = 6'h33 == s2_idx ? ~s2_way[0] : plru1_51; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_345 = 6'h34 == s2_idx ? ~s2_way[0] : plru1_52; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_346 = 6'h35 == s2_idx ? ~s2_way[0] : plru1_53; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_347 = 6'h36 == s2_idx ? ~s2_way[0] : plru1_54; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_348 = 6'h37 == s2_idx ? ~s2_way[0] : plru1_55; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_349 = 6'h38 == s2_idx ? ~s2_way[0] : plru1_56; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_350 = 6'h39 == s2_idx ? ~s2_way[0] : plru1_57; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_351 = 6'h3a == s2_idx ? ~s2_way[0] : plru1_58; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_352 = 6'h3b == s2_idx ? ~s2_way[0] : plru1_59; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_353 = 6'h3c == s2_idx ? ~s2_way[0] : plru1_60; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_354 = 6'h3d == s2_idx ? ~s2_way[0] : plru1_61; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_355 = 6'h3e == s2_idx ? ~s2_way[0] : plru1_62; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_356 = 6'h3f == s2_idx ? ~s2_way[0] : plru1_63; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_357 = 6'h0 == s2_idx ? _plru1_T_1 : plru2_0; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_358 = 6'h1 == s2_idx ? _plru1_T_1 : plru2_1; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_359 = 6'h2 == s2_idx ? _plru1_T_1 : plru2_2; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_360 = 6'h3 == s2_idx ? _plru1_T_1 : plru2_3; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_361 = 6'h4 == s2_idx ? _plru1_T_1 : plru2_4; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_362 = 6'h5 == s2_idx ? _plru1_T_1 : plru2_5; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_363 = 6'h6 == s2_idx ? _plru1_T_1 : plru2_6; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_364 = 6'h7 == s2_idx ? _plru1_T_1 : plru2_7; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_365 = 6'h8 == s2_idx ? _plru1_T_1 : plru2_8; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_366 = 6'h9 == s2_idx ? _plru1_T_1 : plru2_9; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_367 = 6'ha == s2_idx ? _plru1_T_1 : plru2_10; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_368 = 6'hb == s2_idx ? _plru1_T_1 : plru2_11; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_369 = 6'hc == s2_idx ? _plru1_T_1 : plru2_12; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_370 = 6'hd == s2_idx ? _plru1_T_1 : plru2_13; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_371 = 6'he == s2_idx ? _plru1_T_1 : plru2_14; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_372 = 6'hf == s2_idx ? _plru1_T_1 : plru2_15; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_373 = 6'h10 == s2_idx ? _plru1_T_1 : plru2_16; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_374 = 6'h11 == s2_idx ? _plru1_T_1 : plru2_17; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_375 = 6'h12 == s2_idx ? _plru1_T_1 : plru2_18; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_376 = 6'h13 == s2_idx ? _plru1_T_1 : plru2_19; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_377 = 6'h14 == s2_idx ? _plru1_T_1 : plru2_20; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_378 = 6'h15 == s2_idx ? _plru1_T_1 : plru2_21; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_379 = 6'h16 == s2_idx ? _plru1_T_1 : plru2_22; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_380 = 6'h17 == s2_idx ? _plru1_T_1 : plru2_23; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_381 = 6'h18 == s2_idx ? _plru1_T_1 : plru2_24; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_382 = 6'h19 == s2_idx ? _plru1_T_1 : plru2_25; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_383 = 6'h1a == s2_idx ? _plru1_T_1 : plru2_26; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_384 = 6'h1b == s2_idx ? _plru1_T_1 : plru2_27; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_385 = 6'h1c == s2_idx ? _plru1_T_1 : plru2_28; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_386 = 6'h1d == s2_idx ? _plru1_T_1 : plru2_29; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_387 = 6'h1e == s2_idx ? _plru1_T_1 : plru2_30; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_388 = 6'h1f == s2_idx ? _plru1_T_1 : plru2_31; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_389 = 6'h20 == s2_idx ? _plru1_T_1 : plru2_32; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_390 = 6'h21 == s2_idx ? _plru1_T_1 : plru2_33; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_391 = 6'h22 == s2_idx ? _plru1_T_1 : plru2_34; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_392 = 6'h23 == s2_idx ? _plru1_T_1 : plru2_35; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_393 = 6'h24 == s2_idx ? _plru1_T_1 : plru2_36; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_394 = 6'h25 == s2_idx ? _plru1_T_1 : plru2_37; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_395 = 6'h26 == s2_idx ? _plru1_T_1 : plru2_38; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_396 = 6'h27 == s2_idx ? _plru1_T_1 : plru2_39; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_397 = 6'h28 == s2_idx ? _plru1_T_1 : plru2_40; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_398 = 6'h29 == s2_idx ? _plru1_T_1 : plru2_41; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_399 = 6'h2a == s2_idx ? _plru1_T_1 : plru2_42; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_400 = 6'h2b == s2_idx ? _plru1_T_1 : plru2_43; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_401 = 6'h2c == s2_idx ? _plru1_T_1 : plru2_44; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_402 = 6'h2d == s2_idx ? _plru1_T_1 : plru2_45; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_403 = 6'h2e == s2_idx ? _plru1_T_1 : plru2_46; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_404 = 6'h2f == s2_idx ? _plru1_T_1 : plru2_47; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_405 = 6'h30 == s2_idx ? _plru1_T_1 : plru2_48; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_406 = 6'h31 == s2_idx ? _plru1_T_1 : plru2_49; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_407 = 6'h32 == s2_idx ? _plru1_T_1 : plru2_50; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_408 = 6'h33 == s2_idx ? _plru1_T_1 : plru2_51; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_409 = 6'h34 == s2_idx ? _plru1_T_1 : plru2_52; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_410 = 6'h35 == s2_idx ? _plru1_T_1 : plru2_53; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_411 = 6'h36 == s2_idx ? _plru1_T_1 : plru2_54; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_412 = 6'h37 == s2_idx ? _plru1_T_1 : plru2_55; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_413 = 6'h38 == s2_idx ? _plru1_T_1 : plru2_56; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_414 = 6'h39 == s2_idx ? _plru1_T_1 : plru2_57; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_415 = 6'h3a == s2_idx ? _plru1_T_1 : plru2_58; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_416 = 6'h3b == s2_idx ? _plru1_T_1 : plru2_59; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_417 = 6'h3c == s2_idx ? _plru1_T_1 : plru2_60; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_418 = 6'h3d == s2_idx ? _plru1_T_1 : plru2_61; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_419 = 6'h3e == s2_idx ? _plru1_T_1 : plru2_62; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_420 = 6'h3f == s2_idx ? _plru1_T_1 : plru2_63; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_421 = _plru0_T_1 ? _GEN_293 : plru1_0; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_422 = _plru0_T_1 ? _GEN_294 : plru1_1; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_423 = _plru0_T_1 ? _GEN_295 : plru1_2; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_424 = _plru0_T_1 ? _GEN_296 : plru1_3; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_425 = _plru0_T_1 ? _GEN_297 : plru1_4; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_426 = _plru0_T_1 ? _GEN_298 : plru1_5; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_427 = _plru0_T_1 ? _GEN_299 : plru1_6; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_428 = _plru0_T_1 ? _GEN_300 : plru1_7; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_429 = _plru0_T_1 ? _GEN_301 : plru1_8; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_430 = _plru0_T_1 ? _GEN_302 : plru1_9; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_431 = _plru0_T_1 ? _GEN_303 : plru1_10; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_432 = _plru0_T_1 ? _GEN_304 : plru1_11; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_433 = _plru0_T_1 ? _GEN_305 : plru1_12; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_434 = _plru0_T_1 ? _GEN_306 : plru1_13; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_435 = _plru0_T_1 ? _GEN_307 : plru1_14; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_436 = _plru0_T_1 ? _GEN_308 : plru1_15; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_437 = _plru0_T_1 ? _GEN_309 : plru1_16; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_438 = _plru0_T_1 ? _GEN_310 : plru1_17; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_439 = _plru0_T_1 ? _GEN_311 : plru1_18; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_440 = _plru0_T_1 ? _GEN_312 : plru1_19; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_441 = _plru0_T_1 ? _GEN_313 : plru1_20; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_442 = _plru0_T_1 ? _GEN_314 : plru1_21; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_443 = _plru0_T_1 ? _GEN_315 : plru1_22; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_444 = _plru0_T_1 ? _GEN_316 : plru1_23; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_445 = _plru0_T_1 ? _GEN_317 : plru1_24; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_446 = _plru0_T_1 ? _GEN_318 : plru1_25; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_447 = _plru0_T_1 ? _GEN_319 : plru1_26; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_448 = _plru0_T_1 ? _GEN_320 : plru1_27; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_449 = _plru0_T_1 ? _GEN_321 : plru1_28; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_450 = _plru0_T_1 ? _GEN_322 : plru1_29; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_451 = _plru0_T_1 ? _GEN_323 : plru1_30; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_452 = _plru0_T_1 ? _GEN_324 : plru1_31; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_453 = _plru0_T_1 ? _GEN_325 : plru1_32; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_454 = _plru0_T_1 ? _GEN_326 : plru1_33; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_455 = _plru0_T_1 ? _GEN_327 : plru1_34; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_456 = _plru0_T_1 ? _GEN_328 : plru1_35; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_457 = _plru0_T_1 ? _GEN_329 : plru1_36; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_458 = _plru0_T_1 ? _GEN_330 : plru1_37; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_459 = _plru0_T_1 ? _GEN_331 : plru1_38; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_460 = _plru0_T_1 ? _GEN_332 : plru1_39; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_461 = _plru0_T_1 ? _GEN_333 : plru1_40; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_462 = _plru0_T_1 ? _GEN_334 : plru1_41; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_463 = _plru0_T_1 ? _GEN_335 : plru1_42; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_464 = _plru0_T_1 ? _GEN_336 : plru1_43; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_465 = _plru0_T_1 ? _GEN_337 : plru1_44; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_466 = _plru0_T_1 ? _GEN_338 : plru1_45; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_467 = _plru0_T_1 ? _GEN_339 : plru1_46; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_468 = _plru0_T_1 ? _GEN_340 : plru1_47; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_469 = _plru0_T_1 ? _GEN_341 : plru1_48; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_470 = _plru0_T_1 ? _GEN_342 : plru1_49; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_471 = _plru0_T_1 ? _GEN_343 : plru1_50; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_472 = _plru0_T_1 ? _GEN_344 : plru1_51; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_473 = _plru0_T_1 ? _GEN_345 : plru1_52; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_474 = _plru0_T_1 ? _GEN_346 : plru1_53; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_475 = _plru0_T_1 ? _GEN_347 : plru1_54; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_476 = _plru0_T_1 ? _GEN_348 : plru1_55; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_477 = _plru0_T_1 ? _GEN_349 : plru1_56; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_478 = _plru0_T_1 ? _GEN_350 : plru1_57; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_479 = _plru0_T_1 ? _GEN_351 : plru1_58; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_480 = _plru0_T_1 ? _GEN_352 : plru1_59; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_481 = _plru0_T_1 ? _GEN_353 : plru1_60; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_482 = _plru0_T_1 ? _GEN_354 : plru1_61; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_483 = _plru0_T_1 ? _GEN_355 : plru1_62; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_484 = _plru0_T_1 ? _GEN_356 : plru1_63; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_485 = _plru0_T_1 ? plru2_0 : _GEN_357; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_486 = _plru0_T_1 ? plru2_1 : _GEN_358; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_487 = _plru0_T_1 ? plru2_2 : _GEN_359; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_488 = _plru0_T_1 ? plru2_3 : _GEN_360; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_489 = _plru0_T_1 ? plru2_4 : _GEN_361; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_490 = _plru0_T_1 ? plru2_5 : _GEN_362; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_491 = _plru0_T_1 ? plru2_6 : _GEN_363; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_492 = _plru0_T_1 ? plru2_7 : _GEN_364; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_493 = _plru0_T_1 ? plru2_8 : _GEN_365; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_494 = _plru0_T_1 ? plru2_9 : _GEN_366; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_495 = _plru0_T_1 ? plru2_10 : _GEN_367; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_496 = _plru0_T_1 ? plru2_11 : _GEN_368; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_497 = _plru0_T_1 ? plru2_12 : _GEN_369; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_498 = _plru0_T_1 ? plru2_13 : _GEN_370; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_499 = _plru0_T_1 ? plru2_14 : _GEN_371; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_500 = _plru0_T_1 ? plru2_15 : _GEN_372; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_501 = _plru0_T_1 ? plru2_16 : _GEN_373; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_502 = _plru0_T_1 ? plru2_17 : _GEN_374; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_503 = _plru0_T_1 ? plru2_18 : _GEN_375; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_504 = _plru0_T_1 ? plru2_19 : _GEN_376; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_505 = _plru0_T_1 ? plru2_20 : _GEN_377; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_506 = _plru0_T_1 ? plru2_21 : _GEN_378; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_507 = _plru0_T_1 ? plru2_22 : _GEN_379; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_508 = _plru0_T_1 ? plru2_23 : _GEN_380; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_509 = _plru0_T_1 ? plru2_24 : _GEN_381; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_510 = _plru0_T_1 ? plru2_25 : _GEN_382; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_511 = _plru0_T_1 ? plru2_26 : _GEN_383; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_512 = _plru0_T_1 ? plru2_27 : _GEN_384; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_513 = _plru0_T_1 ? plru2_28 : _GEN_385; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_514 = _plru0_T_1 ? plru2_29 : _GEN_386; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_515 = _plru0_T_1 ? plru2_30 : _GEN_387; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_516 = _plru0_T_1 ? plru2_31 : _GEN_388; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_517 = _plru0_T_1 ? plru2_32 : _GEN_389; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_518 = _plru0_T_1 ? plru2_33 : _GEN_390; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_519 = _plru0_T_1 ? plru2_34 : _GEN_391; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_520 = _plru0_T_1 ? plru2_35 : _GEN_392; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_521 = _plru0_T_1 ? plru2_36 : _GEN_393; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_522 = _plru0_T_1 ? plru2_37 : _GEN_394; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_523 = _plru0_T_1 ? plru2_38 : _GEN_395; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_524 = _plru0_T_1 ? plru2_39 : _GEN_396; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_525 = _plru0_T_1 ? plru2_40 : _GEN_397; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_526 = _plru0_T_1 ? plru2_41 : _GEN_398; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_527 = _plru0_T_1 ? plru2_42 : _GEN_399; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_528 = _plru0_T_1 ? plru2_43 : _GEN_400; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_529 = _plru0_T_1 ? plru2_44 : _GEN_401; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_530 = _plru0_T_1 ? plru2_45 : _GEN_402; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_531 = _plru0_T_1 ? plru2_46 : _GEN_403; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_532 = _plru0_T_1 ? plru2_47 : _GEN_404; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_533 = _plru0_T_1 ? plru2_48 : _GEN_405; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_534 = _plru0_T_1 ? plru2_49 : _GEN_406; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_535 = _plru0_T_1 ? plru2_50 : _GEN_407; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_536 = _plru0_T_1 ? plru2_51 : _GEN_408; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_537 = _plru0_T_1 ? plru2_52 : _GEN_409; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_538 = _plru0_T_1 ? plru2_53 : _GEN_410; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_539 = _plru0_T_1 ? plru2_54 : _GEN_411; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_540 = _plru0_T_1 ? plru2_55 : _GEN_412; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_541 = _plru0_T_1 ? plru2_56 : _GEN_413; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_542 = _plru0_T_1 ? plru2_57 : _GEN_414; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_543 = _plru0_T_1 ? plru2_58 : _GEN_415; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_544 = _plru0_T_1 ? plru2_59 : _GEN_416; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_545 = _plru0_T_1 ? plru2_60 : _GEN_417; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_546 = _plru0_T_1 ? plru2_61 : _GEN_418; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_547 = _plru0_T_1 ? plru2_62 : _GEN_419; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_548 = _plru0_T_1 ? plru2_63 : _GEN_420; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _T_6 = s2_way == 2'h0; // @[Cache.scala 295:26]
  wire [7:0] sram_0_io_wdata_lo_lo_lo = s2_wmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] sram_0_io_wdata_lo_lo_hi = s2_wmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] sram_0_io_wdata_lo_hi_lo = s2_wmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] sram_0_io_wdata_lo_hi_hi = s2_wmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] sram_0_io_wdata_hi_lo_lo = s2_wmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] sram_0_io_wdata_hi_lo_hi = s2_wmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] sram_0_io_wdata_hi_hi_lo = s2_wmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] sram_0_io_wdata_hi_hi_hi = s2_wmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _sram_0_io_wdata_T_18 = {sram_0_io_wdata_hi_hi_hi,sram_0_io_wdata_hi_hi_lo,sram_0_io_wdata_hi_lo_hi,
    sram_0_io_wdata_hi_lo_lo,sram_0_io_wdata_lo_hi_hi,sram_0_io_wdata_lo_hi_lo,sram_0_io_wdata_lo_lo_hi,
    sram_0_io_wdata_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] _sram_0_io_wdata_T_19 = s2_wdata & _sram_0_io_wdata_T_18; // @[ID.scala 8:15]
  wire [63:0] _sram_0_io_wdata_T_20 = ~_sram_0_io_wdata_T_18; // @[ID.scala 8:37]
  wire [63:0] _sram_0_io_wdata_T_21 = _GEN_7[127:64] & _sram_0_io_wdata_T_20; // @[ID.scala 8:35]
  wire [63:0] sram_0_io_wdata_hi_1 = _sram_0_io_wdata_T_19 | _sram_0_io_wdata_T_21; // @[ID.scala 8:23]
  wire [127:0] _sram_0_io_wdata_T_22 = {sram_0_io_wdata_hi_1,_GEN_7[63:0]}; // @[Cat.scala 30:58]
  wire [63:0] _sram_0_io_wdata_T_43 = _GEN_7[63:0] & _sram_0_io_wdata_T_20; // @[ID.scala 8:35]
  wire [63:0] sram_0_io_wdata_lo_3 = _sram_0_io_wdata_T_19 | _sram_0_io_wdata_T_43; // @[ID.scala 8:23]
  wire [127:0] _sram_0_io_wdata_T_44 = {_GEN_7[127:64],sram_0_io_wdata_lo_3}; // @[Cat.scala 30:58]
  wire [127:0] _sram_0_io_wdata_T_45 = s2_offs ? _sram_0_io_wdata_T_22 : _sram_0_io_wdata_T_44; // @[Cache.scala 299:38]
  wire  _GEN_741 = s2_way == 2'h0 | fi_ready; // @[Cache.scala 295:35 Cache.scala 296:29]
  wire [5:0] _GEN_743 = s2_way == 2'h0 ? s2_idx : _GEN_3; // @[Cache.scala 295:35 Cache.scala 298:31]
  wire [127:0] _GEN_744 = s2_way == 2'h0 ? _sram_0_io_wdata_T_45 : 128'h0; // @[Cache.scala 295:35 Cache.scala 299:32 Cache.scala 112:16]
  wire  _T_7 = s2_way == 2'h1; // @[Cache.scala 295:26]
  wire  _GEN_745 = s2_way == 2'h1 | fi_ready; // @[Cache.scala 295:35 Cache.scala 296:29]
  wire [5:0] _GEN_747 = s2_way == 2'h1 ? s2_idx : _GEN_3; // @[Cache.scala 295:35 Cache.scala 298:31]
  wire [127:0] _GEN_748 = s2_way == 2'h1 ? _sram_0_io_wdata_T_45 : 128'h0; // @[Cache.scala 295:35 Cache.scala 299:32 Cache.scala 112:16]
  wire  _T_8 = s2_way == 2'h2; // @[Cache.scala 295:26]
  wire  _GEN_749 = s2_way == 2'h2 | fi_ready; // @[Cache.scala 295:35 Cache.scala 296:29]
  wire [5:0] _GEN_751 = s2_way == 2'h2 ? s2_idx : _GEN_3; // @[Cache.scala 295:35 Cache.scala 298:31]
  wire [127:0] _GEN_752 = s2_way == 2'h2 ? _sram_0_io_wdata_T_45 : 128'h0; // @[Cache.scala 295:35 Cache.scala 299:32 Cache.scala 112:16]
  wire  _T_9 = s2_way == 2'h3; // @[Cache.scala 295:26]
  wire  _GEN_753 = s2_way == 2'h3 | fi_ready; // @[Cache.scala 295:35 Cache.scala 296:29]
  wire [5:0] _GEN_755 = s2_way == 2'h3 ? s2_idx : _GEN_3; // @[Cache.scala 295:35 Cache.scala 298:31]
  wire [127:0] _GEN_756 = s2_way == 2'h3 ? _sram_0_io_wdata_T_45 : 128'h0; // @[Cache.scala 295:35 Cache.scala 299:32 Cache.scala 112:16]
  wire [3:0] _GEN_757 = ~s2_hit ? 4'h1 : state; // @[Cache.scala 308:31 Cache.scala 309:17 Cache.scala 207:22]
  wire  _GEN_758 = s2_hit & s2_wen ? _GEN_741 : fi_ready; // @[Cache.scala 293:33]
  wire  _GEN_759 = s2_hit & s2_wen & _T_6; // @[Cache.scala 293:33 Cache.scala 110:14]
  wire [5:0] _GEN_760 = s2_hit & s2_wen ? _GEN_743 : _GEN_3; // @[Cache.scala 293:33]
  wire [127:0] _GEN_761 = s2_hit & s2_wen ? _GEN_744 : 128'h0; // @[Cache.scala 293:33 Cache.scala 112:16]
  wire  _GEN_762 = s2_hit & s2_wen ? _GEN_745 : fi_ready; // @[Cache.scala 293:33]
  wire  _GEN_763 = s2_hit & s2_wen & _T_7; // @[Cache.scala 293:33 Cache.scala 110:14]
  wire [5:0] _GEN_764 = s2_hit & s2_wen ? _GEN_747 : _GEN_3; // @[Cache.scala 293:33]
  wire [127:0] _GEN_765 = s2_hit & s2_wen ? _GEN_748 : 128'h0; // @[Cache.scala 293:33 Cache.scala 112:16]
  wire  _GEN_766 = s2_hit & s2_wen ? _GEN_749 : fi_ready; // @[Cache.scala 293:33]
  wire  _GEN_767 = s2_hit & s2_wen & _T_8; // @[Cache.scala 293:33 Cache.scala 110:14]
  wire [5:0] _GEN_768 = s2_hit & s2_wen ? _GEN_751 : _GEN_3; // @[Cache.scala 293:33]
  wire [127:0] _GEN_769 = s2_hit & s2_wen ? _GEN_752 : 128'h0; // @[Cache.scala 293:33 Cache.scala 112:16]
  wire  _GEN_770 = s2_hit & s2_wen ? _GEN_753 : fi_ready; // @[Cache.scala 293:33]
  wire  _GEN_771 = s2_hit & s2_wen & _T_9; // @[Cache.scala 293:33 Cache.scala 110:14]
  wire [5:0] _GEN_772 = s2_hit & s2_wen ? _GEN_755 : _GEN_3; // @[Cache.scala 293:33]
  wire [127:0] _GEN_773 = s2_hit & s2_wen ? _GEN_756 : 128'h0; // @[Cache.scala 293:33 Cache.scala 112:16]
  wire [3:0] _GEN_774 = s2_hit & s2_wen ? 4'h7 : _GEN_757; // @[Cache.scala 293:33 Cache.scala 307:17]
  wire  _GEN_967 = REG_2 ? _GEN_758 : fi_ready; // @[Cache.scala 289:37]
  wire  _GEN_968 = REG_2 & _GEN_759; // @[Cache.scala 289:37 Cache.scala 110:14]
  wire [5:0] _GEN_969 = REG_2 ? _GEN_760 : _GEN_3; // @[Cache.scala 289:37]
  wire [127:0] _GEN_970 = REG_2 ? _GEN_761 : 128'h0; // @[Cache.scala 289:37 Cache.scala 112:16]
  wire  _GEN_971 = REG_2 ? _GEN_762 : fi_ready; // @[Cache.scala 289:37]
  wire  _GEN_972 = REG_2 & _GEN_763; // @[Cache.scala 289:37 Cache.scala 110:14]
  wire [5:0] _GEN_973 = REG_2 ? _GEN_764 : _GEN_3; // @[Cache.scala 289:37]
  wire [127:0] _GEN_974 = REG_2 ? _GEN_765 : 128'h0; // @[Cache.scala 289:37 Cache.scala 112:16]
  wire  _GEN_975 = REG_2 ? _GEN_766 : fi_ready; // @[Cache.scala 289:37]
  wire  _GEN_976 = REG_2 & _GEN_767; // @[Cache.scala 289:37 Cache.scala 110:14]
  wire [5:0] _GEN_977 = REG_2 ? _GEN_768 : _GEN_3; // @[Cache.scala 289:37]
  wire [127:0] _GEN_978 = REG_2 ? _GEN_769 : 128'h0; // @[Cache.scala 289:37 Cache.scala 112:16]
  wire  _GEN_979 = REG_2 ? _GEN_770 : fi_ready; // @[Cache.scala 289:37]
  wire  _GEN_980 = REG_2 & _GEN_771; // @[Cache.scala 289:37 Cache.scala 110:14]
  wire [5:0] _GEN_981 = REG_2 ? _GEN_772 : _GEN_3; // @[Cache.scala 289:37]
  wire [127:0] _GEN_982 = REG_2 ? _GEN_773 : 128'h0; // @[Cache.scala 289:37 Cache.scala 112:16]
  wire [3:0] _GEN_983 = REG_2 ? _GEN_774 : state; // @[Cache.scala 289:37 Cache.scala 207:22]
  wire  _T_11 = 4'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_984 = _T_12 ? 4'h2 : state; // @[Cache.scala 314:29 Cache.scala 315:15 Cache.scala 207:22]
  wire  _T_13 = 4'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_14 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_985 = ~io_out_resp_bits_rlast ? io_out_resp_bits_rdata : wdata1; // @[Cache.scala 320:37 Cache.scala 321:18 Cache.scala 258:23]
  wire [63:0] _GEN_986 = ~io_out_resp_bits_rlast ? wdata2 : io_out_resp_bits_rdata; // @[Cache.scala 320:37 Cache.scala 259:23 Cache.scala 323:18]
  wire [3:0] _GEN_987 = ~io_out_resp_bits_rlast ? state : 4'h3; // @[Cache.scala 320:37 Cache.scala 207:22 Cache.scala 324:17]
  wire [63:0] _GEN_988 = _T_14 ? _GEN_985 : wdata1; // @[Cache.scala 319:30 Cache.scala 258:23]
  wire [63:0] _GEN_989 = _T_14 ? _GEN_986 : wdata2; // @[Cache.scala 319:30 Cache.scala 259:23]
  wire [3:0] _GEN_990 = _T_14 ? _GEN_987 : state; // @[Cache.scala 319:30 Cache.scala 207:22]
  wire  _T_16 = 4'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_17 = replace_way == 2'h0; // @[Cache.scala 330:27]
  wire [63:0] _sram_0_io_wdata_T_66 = wdata2 & _sram_0_io_wdata_T_20; // @[ID.scala 8:35]
  wire [63:0] sram_0_io_wdata_hi_5 = _sram_0_io_wdata_T_19 | _sram_0_io_wdata_T_66; // @[ID.scala 8:23]
  wire [127:0] _sram_0_io_wdata_T_67 = {sram_0_io_wdata_hi_5,wdata1}; // @[Cat.scala 30:58]
  wire [63:0] _sram_0_io_wdata_T_87 = wdata1 & _sram_0_io_wdata_T_20; // @[ID.scala 8:35]
  wire [63:0] sram_0_io_wdata_lo_6 = _sram_0_io_wdata_T_19 | _sram_0_io_wdata_T_87; // @[ID.scala 8:23]
  wire [127:0] _sram_0_io_wdata_T_88 = {wdata2,sram_0_io_wdata_lo_6}; // @[Cat.scala 30:58]
  wire [127:0] _sram_0_io_wdata_T_89 = s2_offs ? _sram_0_io_wdata_T_67 : _sram_0_io_wdata_T_88; // @[Cache.scala 335:36]
  wire [127:0] _sram_0_io_wdata_T_90 = {wdata2,wdata1}; // @[Cat.scala 30:58]
  wire [127:0] _GEN_991 = s2_wen ? _sram_0_io_wdata_T_89 : _sram_0_io_wdata_T_90; // @[Cache.scala 334:25 Cache.scala 335:30 Cache.scala 339:30]
  wire  _GEN_992 = replace_way == 2'h0 | fi_ready; // @[Cache.scala 330:36 Cache.scala 331:25]
  wire [5:0] _GEN_994 = replace_way == 2'h0 ? s2_idx : _GEN_3; // @[Cache.scala 330:36 Cache.scala 333:27]
  wire [127:0] _GEN_995 = replace_way == 2'h0 ? _GEN_991 : 128'h0; // @[Cache.scala 330:36 Cache.scala 112:16]
  wire [20:0] _GEN_996 = replace_way == 2'h0 ? s2_tag : 21'h0; // @[Cache.scala 330:36 Cache.scala 344:28 Cache.scala 116:16]
  wire  _GEN_997 = replace_way == 2'h0 & s2_wen; // @[Cache.scala 330:36 Cache.scala 346:30 Cache.scala 118:18]
  wire  _T_18 = replace_way == 2'h1; // @[Cache.scala 330:27]
  wire  _GEN_999 = replace_way == 2'h1 | fi_ready; // @[Cache.scala 330:36 Cache.scala 331:25]
  wire [5:0] _GEN_1001 = replace_way == 2'h1 ? s2_idx : _GEN_3; // @[Cache.scala 330:36 Cache.scala 333:27]
  wire [127:0] _GEN_1002 = replace_way == 2'h1 ? _GEN_991 : 128'h0; // @[Cache.scala 330:36 Cache.scala 112:16]
  wire [20:0] _GEN_1003 = replace_way == 2'h1 ? s2_tag : 21'h0; // @[Cache.scala 330:36 Cache.scala 344:28 Cache.scala 116:16]
  wire  _GEN_1004 = replace_way == 2'h1 & s2_wen; // @[Cache.scala 330:36 Cache.scala 346:30 Cache.scala 118:18]
  wire  _T_19 = replace_way == 2'h2; // @[Cache.scala 330:27]
  wire  _GEN_1006 = replace_way == 2'h2 | fi_ready; // @[Cache.scala 330:36 Cache.scala 331:25]
  wire [5:0] _GEN_1008 = replace_way == 2'h2 ? s2_idx : _GEN_3; // @[Cache.scala 330:36 Cache.scala 333:27]
  wire [127:0] _GEN_1009 = replace_way == 2'h2 ? _GEN_991 : 128'h0; // @[Cache.scala 330:36 Cache.scala 112:16]
  wire [20:0] _GEN_1010 = replace_way == 2'h2 ? s2_tag : 21'h0; // @[Cache.scala 330:36 Cache.scala 344:28 Cache.scala 116:16]
  wire  _GEN_1011 = replace_way == 2'h2 & s2_wen; // @[Cache.scala 330:36 Cache.scala 346:30 Cache.scala 118:18]
  wire  _T_20 = replace_way == 2'h3; // @[Cache.scala 330:27]
  wire  _GEN_1013 = replace_way == 2'h3 | fi_ready; // @[Cache.scala 330:36 Cache.scala 331:25]
  wire [5:0] _GEN_1015 = replace_way == 2'h3 ? s2_idx : _GEN_3; // @[Cache.scala 330:36 Cache.scala 333:27]
  wire [127:0] _GEN_1016 = replace_way == 2'h3 ? _GEN_991 : 128'h0; // @[Cache.scala 330:36 Cache.scala 112:16]
  wire [20:0] _GEN_1017 = replace_way == 2'h3 ? s2_tag : 21'h0; // @[Cache.scala 330:36 Cache.scala 344:28 Cache.scala 116:16]
  wire  _GEN_1018 = replace_way == 2'h3 & s2_wen; // @[Cache.scala 330:36 Cache.scala 346:30 Cache.scala 118:18]
  wire  _plru0_T_3 = ~replace_way[1]; // @[Cache.scala 138:19]
  wire  _GEN_1019 = 6'h0 == s2_idx ? ~replace_way[1] : plru0_0; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1020 = 6'h1 == s2_idx ? ~replace_way[1] : plru0_1; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1021 = 6'h2 == s2_idx ? ~replace_way[1] : plru0_2; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1022 = 6'h3 == s2_idx ? ~replace_way[1] : plru0_3; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1023 = 6'h4 == s2_idx ? ~replace_way[1] : plru0_4; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1024 = 6'h5 == s2_idx ? ~replace_way[1] : plru0_5; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1025 = 6'h6 == s2_idx ? ~replace_way[1] : plru0_6; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1026 = 6'h7 == s2_idx ? ~replace_way[1] : plru0_7; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1027 = 6'h8 == s2_idx ? ~replace_way[1] : plru0_8; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1028 = 6'h9 == s2_idx ? ~replace_way[1] : plru0_9; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1029 = 6'ha == s2_idx ? ~replace_way[1] : plru0_10; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1030 = 6'hb == s2_idx ? ~replace_way[1] : plru0_11; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1031 = 6'hc == s2_idx ? ~replace_way[1] : plru0_12; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1032 = 6'hd == s2_idx ? ~replace_way[1] : plru0_13; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1033 = 6'he == s2_idx ? ~replace_way[1] : plru0_14; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1034 = 6'hf == s2_idx ? ~replace_way[1] : plru0_15; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1035 = 6'h10 == s2_idx ? ~replace_way[1] : plru0_16; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1036 = 6'h11 == s2_idx ? ~replace_way[1] : plru0_17; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1037 = 6'h12 == s2_idx ? ~replace_way[1] : plru0_18; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1038 = 6'h13 == s2_idx ? ~replace_way[1] : plru0_19; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1039 = 6'h14 == s2_idx ? ~replace_way[1] : plru0_20; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1040 = 6'h15 == s2_idx ? ~replace_way[1] : plru0_21; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1041 = 6'h16 == s2_idx ? ~replace_way[1] : plru0_22; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1042 = 6'h17 == s2_idx ? ~replace_way[1] : plru0_23; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1043 = 6'h18 == s2_idx ? ~replace_way[1] : plru0_24; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1044 = 6'h19 == s2_idx ? ~replace_way[1] : plru0_25; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1045 = 6'h1a == s2_idx ? ~replace_way[1] : plru0_26; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1046 = 6'h1b == s2_idx ? ~replace_way[1] : plru0_27; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1047 = 6'h1c == s2_idx ? ~replace_way[1] : plru0_28; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1048 = 6'h1d == s2_idx ? ~replace_way[1] : plru0_29; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1049 = 6'h1e == s2_idx ? ~replace_way[1] : plru0_30; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1050 = 6'h1f == s2_idx ? ~replace_way[1] : plru0_31; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1051 = 6'h20 == s2_idx ? ~replace_way[1] : plru0_32; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1052 = 6'h21 == s2_idx ? ~replace_way[1] : plru0_33; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1053 = 6'h22 == s2_idx ? ~replace_way[1] : plru0_34; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1054 = 6'h23 == s2_idx ? ~replace_way[1] : plru0_35; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1055 = 6'h24 == s2_idx ? ~replace_way[1] : plru0_36; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1056 = 6'h25 == s2_idx ? ~replace_way[1] : plru0_37; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1057 = 6'h26 == s2_idx ? ~replace_way[1] : plru0_38; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1058 = 6'h27 == s2_idx ? ~replace_way[1] : plru0_39; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1059 = 6'h28 == s2_idx ? ~replace_way[1] : plru0_40; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1060 = 6'h29 == s2_idx ? ~replace_way[1] : plru0_41; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1061 = 6'h2a == s2_idx ? ~replace_way[1] : plru0_42; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1062 = 6'h2b == s2_idx ? ~replace_way[1] : plru0_43; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1063 = 6'h2c == s2_idx ? ~replace_way[1] : plru0_44; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1064 = 6'h2d == s2_idx ? ~replace_way[1] : plru0_45; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1065 = 6'h2e == s2_idx ? ~replace_way[1] : plru0_46; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1066 = 6'h2f == s2_idx ? ~replace_way[1] : plru0_47; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1067 = 6'h30 == s2_idx ? ~replace_way[1] : plru0_48; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1068 = 6'h31 == s2_idx ? ~replace_way[1] : plru0_49; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1069 = 6'h32 == s2_idx ? ~replace_way[1] : plru0_50; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1070 = 6'h33 == s2_idx ? ~replace_way[1] : plru0_51; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1071 = 6'h34 == s2_idx ? ~replace_way[1] : plru0_52; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1072 = 6'h35 == s2_idx ? ~replace_way[1] : plru0_53; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1073 = 6'h36 == s2_idx ? ~replace_way[1] : plru0_54; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1074 = 6'h37 == s2_idx ? ~replace_way[1] : plru0_55; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1075 = 6'h38 == s2_idx ? ~replace_way[1] : plru0_56; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1076 = 6'h39 == s2_idx ? ~replace_way[1] : plru0_57; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1077 = 6'h3a == s2_idx ? ~replace_way[1] : plru0_58; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1078 = 6'h3b == s2_idx ? ~replace_way[1] : plru0_59; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1079 = 6'h3c == s2_idx ? ~replace_way[1] : plru0_60; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1080 = 6'h3d == s2_idx ? ~replace_way[1] : plru0_61; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1081 = 6'h3e == s2_idx ? ~replace_way[1] : plru0_62; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1082 = 6'h3f == s2_idx ? ~replace_way[1] : plru0_63; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _plru1_T_3 = ~replace_way[0]; // @[Cache.scala 140:21]
  wire  _GEN_1083 = 6'h0 == s2_idx ? ~replace_way[0] : plru1_0; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1084 = 6'h1 == s2_idx ? ~replace_way[0] : plru1_1; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1085 = 6'h2 == s2_idx ? ~replace_way[0] : plru1_2; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1086 = 6'h3 == s2_idx ? ~replace_way[0] : plru1_3; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1087 = 6'h4 == s2_idx ? ~replace_way[0] : plru1_4; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1088 = 6'h5 == s2_idx ? ~replace_way[0] : plru1_5; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1089 = 6'h6 == s2_idx ? ~replace_way[0] : plru1_6; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1090 = 6'h7 == s2_idx ? ~replace_way[0] : plru1_7; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1091 = 6'h8 == s2_idx ? ~replace_way[0] : plru1_8; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1092 = 6'h9 == s2_idx ? ~replace_way[0] : plru1_9; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1093 = 6'ha == s2_idx ? ~replace_way[0] : plru1_10; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1094 = 6'hb == s2_idx ? ~replace_way[0] : plru1_11; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1095 = 6'hc == s2_idx ? ~replace_way[0] : plru1_12; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1096 = 6'hd == s2_idx ? ~replace_way[0] : plru1_13; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1097 = 6'he == s2_idx ? ~replace_way[0] : plru1_14; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1098 = 6'hf == s2_idx ? ~replace_way[0] : plru1_15; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1099 = 6'h10 == s2_idx ? ~replace_way[0] : plru1_16; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1100 = 6'h11 == s2_idx ? ~replace_way[0] : plru1_17; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1101 = 6'h12 == s2_idx ? ~replace_way[0] : plru1_18; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1102 = 6'h13 == s2_idx ? ~replace_way[0] : plru1_19; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1103 = 6'h14 == s2_idx ? ~replace_way[0] : plru1_20; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1104 = 6'h15 == s2_idx ? ~replace_way[0] : plru1_21; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1105 = 6'h16 == s2_idx ? ~replace_way[0] : plru1_22; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1106 = 6'h17 == s2_idx ? ~replace_way[0] : plru1_23; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1107 = 6'h18 == s2_idx ? ~replace_way[0] : plru1_24; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1108 = 6'h19 == s2_idx ? ~replace_way[0] : plru1_25; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1109 = 6'h1a == s2_idx ? ~replace_way[0] : plru1_26; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1110 = 6'h1b == s2_idx ? ~replace_way[0] : plru1_27; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1111 = 6'h1c == s2_idx ? ~replace_way[0] : plru1_28; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1112 = 6'h1d == s2_idx ? ~replace_way[0] : plru1_29; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1113 = 6'h1e == s2_idx ? ~replace_way[0] : plru1_30; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1114 = 6'h1f == s2_idx ? ~replace_way[0] : plru1_31; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1115 = 6'h20 == s2_idx ? ~replace_way[0] : plru1_32; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1116 = 6'h21 == s2_idx ? ~replace_way[0] : plru1_33; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1117 = 6'h22 == s2_idx ? ~replace_way[0] : plru1_34; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1118 = 6'h23 == s2_idx ? ~replace_way[0] : plru1_35; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1119 = 6'h24 == s2_idx ? ~replace_way[0] : plru1_36; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1120 = 6'h25 == s2_idx ? ~replace_way[0] : plru1_37; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1121 = 6'h26 == s2_idx ? ~replace_way[0] : plru1_38; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1122 = 6'h27 == s2_idx ? ~replace_way[0] : plru1_39; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1123 = 6'h28 == s2_idx ? ~replace_way[0] : plru1_40; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1124 = 6'h29 == s2_idx ? ~replace_way[0] : plru1_41; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1125 = 6'h2a == s2_idx ? ~replace_way[0] : plru1_42; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1126 = 6'h2b == s2_idx ? ~replace_way[0] : plru1_43; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1127 = 6'h2c == s2_idx ? ~replace_way[0] : plru1_44; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1128 = 6'h2d == s2_idx ? ~replace_way[0] : plru1_45; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1129 = 6'h2e == s2_idx ? ~replace_way[0] : plru1_46; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1130 = 6'h2f == s2_idx ? ~replace_way[0] : plru1_47; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1131 = 6'h30 == s2_idx ? ~replace_way[0] : plru1_48; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1132 = 6'h31 == s2_idx ? ~replace_way[0] : plru1_49; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1133 = 6'h32 == s2_idx ? ~replace_way[0] : plru1_50; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1134 = 6'h33 == s2_idx ? ~replace_way[0] : plru1_51; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1135 = 6'h34 == s2_idx ? ~replace_way[0] : plru1_52; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1136 = 6'h35 == s2_idx ? ~replace_way[0] : plru1_53; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1137 = 6'h36 == s2_idx ? ~replace_way[0] : plru1_54; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1138 = 6'h37 == s2_idx ? ~replace_way[0] : plru1_55; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1139 = 6'h38 == s2_idx ? ~replace_way[0] : plru1_56; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1140 = 6'h39 == s2_idx ? ~replace_way[0] : plru1_57; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1141 = 6'h3a == s2_idx ? ~replace_way[0] : plru1_58; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1142 = 6'h3b == s2_idx ? ~replace_way[0] : plru1_59; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1143 = 6'h3c == s2_idx ? ~replace_way[0] : plru1_60; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1144 = 6'h3d == s2_idx ? ~replace_way[0] : plru1_61; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1145 = 6'h3e == s2_idx ? ~replace_way[0] : plru1_62; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1146 = 6'h3f == s2_idx ? ~replace_way[0] : plru1_63; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1147 = 6'h0 == s2_idx ? _plru1_T_3 : plru2_0; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1148 = 6'h1 == s2_idx ? _plru1_T_3 : plru2_1; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1149 = 6'h2 == s2_idx ? _plru1_T_3 : plru2_2; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1150 = 6'h3 == s2_idx ? _plru1_T_3 : plru2_3; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1151 = 6'h4 == s2_idx ? _plru1_T_3 : plru2_4; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1152 = 6'h5 == s2_idx ? _plru1_T_3 : plru2_5; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1153 = 6'h6 == s2_idx ? _plru1_T_3 : plru2_6; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1154 = 6'h7 == s2_idx ? _plru1_T_3 : plru2_7; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1155 = 6'h8 == s2_idx ? _plru1_T_3 : plru2_8; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1156 = 6'h9 == s2_idx ? _plru1_T_3 : plru2_9; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1157 = 6'ha == s2_idx ? _plru1_T_3 : plru2_10; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1158 = 6'hb == s2_idx ? _plru1_T_3 : plru2_11; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1159 = 6'hc == s2_idx ? _plru1_T_3 : plru2_12; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1160 = 6'hd == s2_idx ? _plru1_T_3 : plru2_13; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1161 = 6'he == s2_idx ? _plru1_T_3 : plru2_14; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1162 = 6'hf == s2_idx ? _plru1_T_3 : plru2_15; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1163 = 6'h10 == s2_idx ? _plru1_T_3 : plru2_16; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1164 = 6'h11 == s2_idx ? _plru1_T_3 : plru2_17; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1165 = 6'h12 == s2_idx ? _plru1_T_3 : plru2_18; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1166 = 6'h13 == s2_idx ? _plru1_T_3 : plru2_19; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1167 = 6'h14 == s2_idx ? _plru1_T_3 : plru2_20; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1168 = 6'h15 == s2_idx ? _plru1_T_3 : plru2_21; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1169 = 6'h16 == s2_idx ? _plru1_T_3 : plru2_22; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1170 = 6'h17 == s2_idx ? _plru1_T_3 : plru2_23; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1171 = 6'h18 == s2_idx ? _plru1_T_3 : plru2_24; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1172 = 6'h19 == s2_idx ? _plru1_T_3 : plru2_25; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1173 = 6'h1a == s2_idx ? _plru1_T_3 : plru2_26; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1174 = 6'h1b == s2_idx ? _plru1_T_3 : plru2_27; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1175 = 6'h1c == s2_idx ? _plru1_T_3 : plru2_28; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1176 = 6'h1d == s2_idx ? _plru1_T_3 : plru2_29; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1177 = 6'h1e == s2_idx ? _plru1_T_3 : plru2_30; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1178 = 6'h1f == s2_idx ? _plru1_T_3 : plru2_31; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1179 = 6'h20 == s2_idx ? _plru1_T_3 : plru2_32; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1180 = 6'h21 == s2_idx ? _plru1_T_3 : plru2_33; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1181 = 6'h22 == s2_idx ? _plru1_T_3 : plru2_34; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1182 = 6'h23 == s2_idx ? _plru1_T_3 : plru2_35; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1183 = 6'h24 == s2_idx ? _plru1_T_3 : plru2_36; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1184 = 6'h25 == s2_idx ? _plru1_T_3 : plru2_37; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1185 = 6'h26 == s2_idx ? _plru1_T_3 : plru2_38; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1186 = 6'h27 == s2_idx ? _plru1_T_3 : plru2_39; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1187 = 6'h28 == s2_idx ? _plru1_T_3 : plru2_40; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1188 = 6'h29 == s2_idx ? _plru1_T_3 : plru2_41; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1189 = 6'h2a == s2_idx ? _plru1_T_3 : plru2_42; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1190 = 6'h2b == s2_idx ? _plru1_T_3 : plru2_43; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1191 = 6'h2c == s2_idx ? _plru1_T_3 : plru2_44; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1192 = 6'h2d == s2_idx ? _plru1_T_3 : plru2_45; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1193 = 6'h2e == s2_idx ? _plru1_T_3 : plru2_46; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1194 = 6'h2f == s2_idx ? _plru1_T_3 : plru2_47; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1195 = 6'h30 == s2_idx ? _plru1_T_3 : plru2_48; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1196 = 6'h31 == s2_idx ? _plru1_T_3 : plru2_49; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1197 = 6'h32 == s2_idx ? _plru1_T_3 : plru2_50; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1198 = 6'h33 == s2_idx ? _plru1_T_3 : plru2_51; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1199 = 6'h34 == s2_idx ? _plru1_T_3 : plru2_52; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1200 = 6'h35 == s2_idx ? _plru1_T_3 : plru2_53; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1201 = 6'h36 == s2_idx ? _plru1_T_3 : plru2_54; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1202 = 6'h37 == s2_idx ? _plru1_T_3 : plru2_55; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1203 = 6'h38 == s2_idx ? _plru1_T_3 : plru2_56; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1204 = 6'h39 == s2_idx ? _plru1_T_3 : plru2_57; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1205 = 6'h3a == s2_idx ? _plru1_T_3 : plru2_58; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1206 = 6'h3b == s2_idx ? _plru1_T_3 : plru2_59; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1207 = 6'h3c == s2_idx ? _plru1_T_3 : plru2_60; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1208 = 6'h3d == s2_idx ? _plru1_T_3 : plru2_61; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1209 = 6'h3e == s2_idx ? _plru1_T_3 : plru2_62; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1210 = 6'h3f == s2_idx ? _plru1_T_3 : plru2_63; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1211 = _plru0_T_3 ? _GEN_1083 : plru1_0; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1212 = _plru0_T_3 ? _GEN_1084 : plru1_1; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1213 = _plru0_T_3 ? _GEN_1085 : plru1_2; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1214 = _plru0_T_3 ? _GEN_1086 : plru1_3; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1215 = _plru0_T_3 ? _GEN_1087 : plru1_4; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1216 = _plru0_T_3 ? _GEN_1088 : plru1_5; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1217 = _plru0_T_3 ? _GEN_1089 : plru1_6; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1218 = _plru0_T_3 ? _GEN_1090 : plru1_7; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1219 = _plru0_T_3 ? _GEN_1091 : plru1_8; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1220 = _plru0_T_3 ? _GEN_1092 : plru1_9; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1221 = _plru0_T_3 ? _GEN_1093 : plru1_10; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1222 = _plru0_T_3 ? _GEN_1094 : plru1_11; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1223 = _plru0_T_3 ? _GEN_1095 : plru1_12; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1224 = _plru0_T_3 ? _GEN_1096 : plru1_13; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1225 = _plru0_T_3 ? _GEN_1097 : plru1_14; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1226 = _plru0_T_3 ? _GEN_1098 : plru1_15; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1227 = _plru0_T_3 ? _GEN_1099 : plru1_16; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1228 = _plru0_T_3 ? _GEN_1100 : plru1_17; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1229 = _plru0_T_3 ? _GEN_1101 : plru1_18; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1230 = _plru0_T_3 ? _GEN_1102 : plru1_19; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1231 = _plru0_T_3 ? _GEN_1103 : plru1_20; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1232 = _plru0_T_3 ? _GEN_1104 : plru1_21; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1233 = _plru0_T_3 ? _GEN_1105 : plru1_22; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1234 = _plru0_T_3 ? _GEN_1106 : plru1_23; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1235 = _plru0_T_3 ? _GEN_1107 : plru1_24; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1236 = _plru0_T_3 ? _GEN_1108 : plru1_25; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1237 = _plru0_T_3 ? _GEN_1109 : plru1_26; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1238 = _plru0_T_3 ? _GEN_1110 : plru1_27; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1239 = _plru0_T_3 ? _GEN_1111 : plru1_28; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1240 = _plru0_T_3 ? _GEN_1112 : plru1_29; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1241 = _plru0_T_3 ? _GEN_1113 : plru1_30; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1242 = _plru0_T_3 ? _GEN_1114 : plru1_31; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1243 = _plru0_T_3 ? _GEN_1115 : plru1_32; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1244 = _plru0_T_3 ? _GEN_1116 : plru1_33; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1245 = _plru0_T_3 ? _GEN_1117 : plru1_34; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1246 = _plru0_T_3 ? _GEN_1118 : plru1_35; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1247 = _plru0_T_3 ? _GEN_1119 : plru1_36; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1248 = _plru0_T_3 ? _GEN_1120 : plru1_37; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1249 = _plru0_T_3 ? _GEN_1121 : plru1_38; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1250 = _plru0_T_3 ? _GEN_1122 : plru1_39; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1251 = _plru0_T_3 ? _GEN_1123 : plru1_40; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1252 = _plru0_T_3 ? _GEN_1124 : plru1_41; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1253 = _plru0_T_3 ? _GEN_1125 : plru1_42; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1254 = _plru0_T_3 ? _GEN_1126 : plru1_43; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1255 = _plru0_T_3 ? _GEN_1127 : plru1_44; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1256 = _plru0_T_3 ? _GEN_1128 : plru1_45; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1257 = _plru0_T_3 ? _GEN_1129 : plru1_46; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1258 = _plru0_T_3 ? _GEN_1130 : plru1_47; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1259 = _plru0_T_3 ? _GEN_1131 : plru1_48; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1260 = _plru0_T_3 ? _GEN_1132 : plru1_49; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1261 = _plru0_T_3 ? _GEN_1133 : plru1_50; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1262 = _plru0_T_3 ? _GEN_1134 : plru1_51; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1263 = _plru0_T_3 ? _GEN_1135 : plru1_52; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1264 = _plru0_T_3 ? _GEN_1136 : plru1_53; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1265 = _plru0_T_3 ? _GEN_1137 : plru1_54; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1266 = _plru0_T_3 ? _GEN_1138 : plru1_55; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1267 = _plru0_T_3 ? _GEN_1139 : plru1_56; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1268 = _plru0_T_3 ? _GEN_1140 : plru1_57; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1269 = _plru0_T_3 ? _GEN_1141 : plru1_58; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1270 = _plru0_T_3 ? _GEN_1142 : plru1_59; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1271 = _plru0_T_3 ? _GEN_1143 : plru1_60; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1272 = _plru0_T_3 ? _GEN_1144 : plru1_61; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1273 = _plru0_T_3 ? _GEN_1145 : plru1_62; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1274 = _plru0_T_3 ? _GEN_1146 : plru1_63; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1275 = _plru0_T_3 ? plru2_0 : _GEN_1147; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1276 = _plru0_T_3 ? plru2_1 : _GEN_1148; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1277 = _plru0_T_3 ? plru2_2 : _GEN_1149; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1278 = _plru0_T_3 ? plru2_3 : _GEN_1150; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1279 = _plru0_T_3 ? plru2_4 : _GEN_1151; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1280 = _plru0_T_3 ? plru2_5 : _GEN_1152; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1281 = _plru0_T_3 ? plru2_6 : _GEN_1153; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1282 = _plru0_T_3 ? plru2_7 : _GEN_1154; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1283 = _plru0_T_3 ? plru2_8 : _GEN_1155; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1284 = _plru0_T_3 ? plru2_9 : _GEN_1156; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1285 = _plru0_T_3 ? plru2_10 : _GEN_1157; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1286 = _plru0_T_3 ? plru2_11 : _GEN_1158; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1287 = _plru0_T_3 ? plru2_12 : _GEN_1159; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1288 = _plru0_T_3 ? plru2_13 : _GEN_1160; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1289 = _plru0_T_3 ? plru2_14 : _GEN_1161; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1290 = _plru0_T_3 ? plru2_15 : _GEN_1162; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1291 = _plru0_T_3 ? plru2_16 : _GEN_1163; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1292 = _plru0_T_3 ? plru2_17 : _GEN_1164; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1293 = _plru0_T_3 ? plru2_18 : _GEN_1165; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1294 = _plru0_T_3 ? plru2_19 : _GEN_1166; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1295 = _plru0_T_3 ? plru2_20 : _GEN_1167; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1296 = _plru0_T_3 ? plru2_21 : _GEN_1168; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1297 = _plru0_T_3 ? plru2_22 : _GEN_1169; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1298 = _plru0_T_3 ? plru2_23 : _GEN_1170; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1299 = _plru0_T_3 ? plru2_24 : _GEN_1171; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1300 = _plru0_T_3 ? plru2_25 : _GEN_1172; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1301 = _plru0_T_3 ? plru2_26 : _GEN_1173; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1302 = _plru0_T_3 ? plru2_27 : _GEN_1174; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1303 = _plru0_T_3 ? plru2_28 : _GEN_1175; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1304 = _plru0_T_3 ? plru2_29 : _GEN_1176; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1305 = _plru0_T_3 ? plru2_30 : _GEN_1177; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1306 = _plru0_T_3 ? plru2_31 : _GEN_1178; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1307 = _plru0_T_3 ? plru2_32 : _GEN_1179; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1308 = _plru0_T_3 ? plru2_33 : _GEN_1180; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1309 = _plru0_T_3 ? plru2_34 : _GEN_1181; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1310 = _plru0_T_3 ? plru2_35 : _GEN_1182; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1311 = _plru0_T_3 ? plru2_36 : _GEN_1183; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1312 = _plru0_T_3 ? plru2_37 : _GEN_1184; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1313 = _plru0_T_3 ? plru2_38 : _GEN_1185; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1314 = _plru0_T_3 ? plru2_39 : _GEN_1186; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1315 = _plru0_T_3 ? plru2_40 : _GEN_1187; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1316 = _plru0_T_3 ? plru2_41 : _GEN_1188; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1317 = _plru0_T_3 ? plru2_42 : _GEN_1189; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1318 = _plru0_T_3 ? plru2_43 : _GEN_1190; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1319 = _plru0_T_3 ? plru2_44 : _GEN_1191; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1320 = _plru0_T_3 ? plru2_45 : _GEN_1192; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1321 = _plru0_T_3 ? plru2_46 : _GEN_1193; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1322 = _plru0_T_3 ? plru2_47 : _GEN_1194; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1323 = _plru0_T_3 ? plru2_48 : _GEN_1195; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1324 = _plru0_T_3 ? plru2_49 : _GEN_1196; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1325 = _plru0_T_3 ? plru2_50 : _GEN_1197; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1326 = _plru0_T_3 ? plru2_51 : _GEN_1198; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1327 = _plru0_T_3 ? plru2_52 : _GEN_1199; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1328 = _plru0_T_3 ? plru2_53 : _GEN_1200; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1329 = _plru0_T_3 ? plru2_54 : _GEN_1201; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1330 = _plru0_T_3 ? plru2_55 : _GEN_1202; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1331 = _plru0_T_3 ? plru2_56 : _GEN_1203; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1332 = _plru0_T_3 ? plru2_57 : _GEN_1204; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1333 = _plru0_T_3 ? plru2_58 : _GEN_1205; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1334 = _plru0_T_3 ? plru2_59 : _GEN_1206; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1335 = _plru0_T_3 ? plru2_60 : _GEN_1207; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1336 = _plru0_T_3 ? plru2_61 : _GEN_1208; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1337 = _plru0_T_3 ? plru2_62 : _GEN_1209; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1338 = _plru0_T_3 ? plru2_63 : _GEN_1210; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire [3:0] _GEN_1339 = s2_reg_dirty ? 4'h4 : 4'h7; // @[Cache.scala 349:27 Cache.scala 350:15 Cache.scala 353:15]
  wire  _GEN_1340 = s2_reg_dirty ? plru0_0 : _GEN_1019; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1341 = s2_reg_dirty ? plru0_1 : _GEN_1020; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1342 = s2_reg_dirty ? plru0_2 : _GEN_1021; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1343 = s2_reg_dirty ? plru0_3 : _GEN_1022; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1344 = s2_reg_dirty ? plru0_4 : _GEN_1023; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1345 = s2_reg_dirty ? plru0_5 : _GEN_1024; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1346 = s2_reg_dirty ? plru0_6 : _GEN_1025; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1347 = s2_reg_dirty ? plru0_7 : _GEN_1026; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1348 = s2_reg_dirty ? plru0_8 : _GEN_1027; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1349 = s2_reg_dirty ? plru0_9 : _GEN_1028; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1350 = s2_reg_dirty ? plru0_10 : _GEN_1029; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1351 = s2_reg_dirty ? plru0_11 : _GEN_1030; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1352 = s2_reg_dirty ? plru0_12 : _GEN_1031; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1353 = s2_reg_dirty ? plru0_13 : _GEN_1032; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1354 = s2_reg_dirty ? plru0_14 : _GEN_1033; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1355 = s2_reg_dirty ? plru0_15 : _GEN_1034; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1356 = s2_reg_dirty ? plru0_16 : _GEN_1035; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1357 = s2_reg_dirty ? plru0_17 : _GEN_1036; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1358 = s2_reg_dirty ? plru0_18 : _GEN_1037; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1359 = s2_reg_dirty ? plru0_19 : _GEN_1038; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1360 = s2_reg_dirty ? plru0_20 : _GEN_1039; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1361 = s2_reg_dirty ? plru0_21 : _GEN_1040; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1362 = s2_reg_dirty ? plru0_22 : _GEN_1041; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1363 = s2_reg_dirty ? plru0_23 : _GEN_1042; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1364 = s2_reg_dirty ? plru0_24 : _GEN_1043; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1365 = s2_reg_dirty ? plru0_25 : _GEN_1044; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1366 = s2_reg_dirty ? plru0_26 : _GEN_1045; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1367 = s2_reg_dirty ? plru0_27 : _GEN_1046; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1368 = s2_reg_dirty ? plru0_28 : _GEN_1047; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1369 = s2_reg_dirty ? plru0_29 : _GEN_1048; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1370 = s2_reg_dirty ? plru0_30 : _GEN_1049; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1371 = s2_reg_dirty ? plru0_31 : _GEN_1050; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1372 = s2_reg_dirty ? plru0_32 : _GEN_1051; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1373 = s2_reg_dirty ? plru0_33 : _GEN_1052; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1374 = s2_reg_dirty ? plru0_34 : _GEN_1053; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1375 = s2_reg_dirty ? plru0_35 : _GEN_1054; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1376 = s2_reg_dirty ? plru0_36 : _GEN_1055; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1377 = s2_reg_dirty ? plru0_37 : _GEN_1056; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1378 = s2_reg_dirty ? plru0_38 : _GEN_1057; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1379 = s2_reg_dirty ? plru0_39 : _GEN_1058; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1380 = s2_reg_dirty ? plru0_40 : _GEN_1059; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1381 = s2_reg_dirty ? plru0_41 : _GEN_1060; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1382 = s2_reg_dirty ? plru0_42 : _GEN_1061; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1383 = s2_reg_dirty ? plru0_43 : _GEN_1062; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1384 = s2_reg_dirty ? plru0_44 : _GEN_1063; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1385 = s2_reg_dirty ? plru0_45 : _GEN_1064; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1386 = s2_reg_dirty ? plru0_46 : _GEN_1065; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1387 = s2_reg_dirty ? plru0_47 : _GEN_1066; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1388 = s2_reg_dirty ? plru0_48 : _GEN_1067; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1389 = s2_reg_dirty ? plru0_49 : _GEN_1068; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1390 = s2_reg_dirty ? plru0_50 : _GEN_1069; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1391 = s2_reg_dirty ? plru0_51 : _GEN_1070; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1392 = s2_reg_dirty ? plru0_52 : _GEN_1071; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1393 = s2_reg_dirty ? plru0_53 : _GEN_1072; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1394 = s2_reg_dirty ? plru0_54 : _GEN_1073; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1395 = s2_reg_dirty ? plru0_55 : _GEN_1074; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1396 = s2_reg_dirty ? plru0_56 : _GEN_1075; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1397 = s2_reg_dirty ? plru0_57 : _GEN_1076; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1398 = s2_reg_dirty ? plru0_58 : _GEN_1077; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1399 = s2_reg_dirty ? plru0_59 : _GEN_1078; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1400 = s2_reg_dirty ? plru0_60 : _GEN_1079; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1401 = s2_reg_dirty ? plru0_61 : _GEN_1080; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1402 = s2_reg_dirty ? plru0_62 : _GEN_1081; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1403 = s2_reg_dirty ? plru0_63 : _GEN_1082; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1404 = s2_reg_dirty ? plru1_0 : _GEN_1211; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1405 = s2_reg_dirty ? plru1_1 : _GEN_1212; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1406 = s2_reg_dirty ? plru1_2 : _GEN_1213; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1407 = s2_reg_dirty ? plru1_3 : _GEN_1214; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1408 = s2_reg_dirty ? plru1_4 : _GEN_1215; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1409 = s2_reg_dirty ? plru1_5 : _GEN_1216; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1410 = s2_reg_dirty ? plru1_6 : _GEN_1217; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1411 = s2_reg_dirty ? plru1_7 : _GEN_1218; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1412 = s2_reg_dirty ? plru1_8 : _GEN_1219; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1413 = s2_reg_dirty ? plru1_9 : _GEN_1220; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1414 = s2_reg_dirty ? plru1_10 : _GEN_1221; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1415 = s2_reg_dirty ? plru1_11 : _GEN_1222; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1416 = s2_reg_dirty ? plru1_12 : _GEN_1223; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1417 = s2_reg_dirty ? plru1_13 : _GEN_1224; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1418 = s2_reg_dirty ? plru1_14 : _GEN_1225; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1419 = s2_reg_dirty ? plru1_15 : _GEN_1226; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1420 = s2_reg_dirty ? plru1_16 : _GEN_1227; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1421 = s2_reg_dirty ? plru1_17 : _GEN_1228; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1422 = s2_reg_dirty ? plru1_18 : _GEN_1229; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1423 = s2_reg_dirty ? plru1_19 : _GEN_1230; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1424 = s2_reg_dirty ? plru1_20 : _GEN_1231; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1425 = s2_reg_dirty ? plru1_21 : _GEN_1232; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1426 = s2_reg_dirty ? plru1_22 : _GEN_1233; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1427 = s2_reg_dirty ? plru1_23 : _GEN_1234; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1428 = s2_reg_dirty ? plru1_24 : _GEN_1235; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1429 = s2_reg_dirty ? plru1_25 : _GEN_1236; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1430 = s2_reg_dirty ? plru1_26 : _GEN_1237; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1431 = s2_reg_dirty ? plru1_27 : _GEN_1238; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1432 = s2_reg_dirty ? plru1_28 : _GEN_1239; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1433 = s2_reg_dirty ? plru1_29 : _GEN_1240; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1434 = s2_reg_dirty ? plru1_30 : _GEN_1241; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1435 = s2_reg_dirty ? plru1_31 : _GEN_1242; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1436 = s2_reg_dirty ? plru1_32 : _GEN_1243; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1437 = s2_reg_dirty ? plru1_33 : _GEN_1244; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1438 = s2_reg_dirty ? plru1_34 : _GEN_1245; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1439 = s2_reg_dirty ? plru1_35 : _GEN_1246; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1440 = s2_reg_dirty ? plru1_36 : _GEN_1247; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1441 = s2_reg_dirty ? plru1_37 : _GEN_1248; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1442 = s2_reg_dirty ? plru1_38 : _GEN_1249; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1443 = s2_reg_dirty ? plru1_39 : _GEN_1250; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1444 = s2_reg_dirty ? plru1_40 : _GEN_1251; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1445 = s2_reg_dirty ? plru1_41 : _GEN_1252; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1446 = s2_reg_dirty ? plru1_42 : _GEN_1253; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1447 = s2_reg_dirty ? plru1_43 : _GEN_1254; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1448 = s2_reg_dirty ? plru1_44 : _GEN_1255; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1449 = s2_reg_dirty ? plru1_45 : _GEN_1256; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1450 = s2_reg_dirty ? plru1_46 : _GEN_1257; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1451 = s2_reg_dirty ? plru1_47 : _GEN_1258; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1452 = s2_reg_dirty ? plru1_48 : _GEN_1259; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1453 = s2_reg_dirty ? plru1_49 : _GEN_1260; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1454 = s2_reg_dirty ? plru1_50 : _GEN_1261; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1455 = s2_reg_dirty ? plru1_51 : _GEN_1262; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1456 = s2_reg_dirty ? plru1_52 : _GEN_1263; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1457 = s2_reg_dirty ? plru1_53 : _GEN_1264; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1458 = s2_reg_dirty ? plru1_54 : _GEN_1265; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1459 = s2_reg_dirty ? plru1_55 : _GEN_1266; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1460 = s2_reg_dirty ? plru1_56 : _GEN_1267; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1461 = s2_reg_dirty ? plru1_57 : _GEN_1268; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1462 = s2_reg_dirty ? plru1_58 : _GEN_1269; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1463 = s2_reg_dirty ? plru1_59 : _GEN_1270; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1464 = s2_reg_dirty ? plru1_60 : _GEN_1271; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1465 = s2_reg_dirty ? plru1_61 : _GEN_1272; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1466 = s2_reg_dirty ? plru1_62 : _GEN_1273; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1467 = s2_reg_dirty ? plru1_63 : _GEN_1274; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1468 = s2_reg_dirty ? plru2_0 : _GEN_1275; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1469 = s2_reg_dirty ? plru2_1 : _GEN_1276; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1470 = s2_reg_dirty ? plru2_2 : _GEN_1277; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1471 = s2_reg_dirty ? plru2_3 : _GEN_1278; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1472 = s2_reg_dirty ? plru2_4 : _GEN_1279; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1473 = s2_reg_dirty ? plru2_5 : _GEN_1280; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1474 = s2_reg_dirty ? plru2_6 : _GEN_1281; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1475 = s2_reg_dirty ? plru2_7 : _GEN_1282; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1476 = s2_reg_dirty ? plru2_8 : _GEN_1283; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1477 = s2_reg_dirty ? plru2_9 : _GEN_1284; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1478 = s2_reg_dirty ? plru2_10 : _GEN_1285; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1479 = s2_reg_dirty ? plru2_11 : _GEN_1286; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1480 = s2_reg_dirty ? plru2_12 : _GEN_1287; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1481 = s2_reg_dirty ? plru2_13 : _GEN_1288; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1482 = s2_reg_dirty ? plru2_14 : _GEN_1289; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1483 = s2_reg_dirty ? plru2_15 : _GEN_1290; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1484 = s2_reg_dirty ? plru2_16 : _GEN_1291; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1485 = s2_reg_dirty ? plru2_17 : _GEN_1292; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1486 = s2_reg_dirty ? plru2_18 : _GEN_1293; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1487 = s2_reg_dirty ? plru2_19 : _GEN_1294; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1488 = s2_reg_dirty ? plru2_20 : _GEN_1295; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1489 = s2_reg_dirty ? plru2_21 : _GEN_1296; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1490 = s2_reg_dirty ? plru2_22 : _GEN_1297; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1491 = s2_reg_dirty ? plru2_23 : _GEN_1298; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1492 = s2_reg_dirty ? plru2_24 : _GEN_1299; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1493 = s2_reg_dirty ? plru2_25 : _GEN_1300; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1494 = s2_reg_dirty ? plru2_26 : _GEN_1301; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1495 = s2_reg_dirty ? plru2_27 : _GEN_1302; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1496 = s2_reg_dirty ? plru2_28 : _GEN_1303; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1497 = s2_reg_dirty ? plru2_29 : _GEN_1304; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1498 = s2_reg_dirty ? plru2_30 : _GEN_1305; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1499 = s2_reg_dirty ? plru2_31 : _GEN_1306; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1500 = s2_reg_dirty ? plru2_32 : _GEN_1307; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1501 = s2_reg_dirty ? plru2_33 : _GEN_1308; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1502 = s2_reg_dirty ? plru2_34 : _GEN_1309; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1503 = s2_reg_dirty ? plru2_35 : _GEN_1310; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1504 = s2_reg_dirty ? plru2_36 : _GEN_1311; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1505 = s2_reg_dirty ? plru2_37 : _GEN_1312; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1506 = s2_reg_dirty ? plru2_38 : _GEN_1313; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1507 = s2_reg_dirty ? plru2_39 : _GEN_1314; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1508 = s2_reg_dirty ? plru2_40 : _GEN_1315; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1509 = s2_reg_dirty ? plru2_41 : _GEN_1316; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1510 = s2_reg_dirty ? plru2_42 : _GEN_1317; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1511 = s2_reg_dirty ? plru2_43 : _GEN_1318; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1512 = s2_reg_dirty ? plru2_44 : _GEN_1319; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1513 = s2_reg_dirty ? plru2_45 : _GEN_1320; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1514 = s2_reg_dirty ? plru2_46 : _GEN_1321; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1515 = s2_reg_dirty ? plru2_47 : _GEN_1322; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1516 = s2_reg_dirty ? plru2_48 : _GEN_1323; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1517 = s2_reg_dirty ? plru2_49 : _GEN_1324; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1518 = s2_reg_dirty ? plru2_50 : _GEN_1325; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1519 = s2_reg_dirty ? plru2_51 : _GEN_1326; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1520 = s2_reg_dirty ? plru2_52 : _GEN_1327; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1521 = s2_reg_dirty ? plru2_53 : _GEN_1328; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1522 = s2_reg_dirty ? plru2_54 : _GEN_1329; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1523 = s2_reg_dirty ? plru2_55 : _GEN_1330; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1524 = s2_reg_dirty ? plru2_56 : _GEN_1331; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1525 = s2_reg_dirty ? plru2_57 : _GEN_1332; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1526 = s2_reg_dirty ? plru2_58 : _GEN_1333; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1527 = s2_reg_dirty ? plru2_59 : _GEN_1334; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1528 = s2_reg_dirty ? plru2_60 : _GEN_1335; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1529 = s2_reg_dirty ? plru2_61 : _GEN_1336; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1530 = s2_reg_dirty ? plru2_62 : _GEN_1337; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1531 = s2_reg_dirty ? plru2_63 : _GEN_1338; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _T_23 = 4'h4 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_1532 = _T_12 ? 4'h5 : state; // @[Cache.scala 357:29 Cache.scala 358:15 Cache.scala 207:22]
  wire  _T_25 = 4'h5 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_1533 = _T_12 ? 4'h6 : state; // @[Cache.scala 362:29 Cache.scala 363:15 Cache.scala 207:22]
  wire  _T_27 = 4'h6 == state; // @[Conditional.scala 37:30]
  wire  _GEN_1854 = _T_14 ? _GEN_1019 : plru0_0; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1855 = _T_14 ? _GEN_1020 : plru0_1; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1856 = _T_14 ? _GEN_1021 : plru0_2; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1857 = _T_14 ? _GEN_1022 : plru0_3; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1858 = _T_14 ? _GEN_1023 : plru0_4; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1859 = _T_14 ? _GEN_1024 : plru0_5; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1860 = _T_14 ? _GEN_1025 : plru0_6; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1861 = _T_14 ? _GEN_1026 : plru0_7; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1862 = _T_14 ? _GEN_1027 : plru0_8; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1863 = _T_14 ? _GEN_1028 : plru0_9; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1864 = _T_14 ? _GEN_1029 : plru0_10; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1865 = _T_14 ? _GEN_1030 : plru0_11; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1866 = _T_14 ? _GEN_1031 : plru0_12; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1867 = _T_14 ? _GEN_1032 : plru0_13; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1868 = _T_14 ? _GEN_1033 : plru0_14; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1869 = _T_14 ? _GEN_1034 : plru0_15; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1870 = _T_14 ? _GEN_1035 : plru0_16; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1871 = _T_14 ? _GEN_1036 : plru0_17; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1872 = _T_14 ? _GEN_1037 : plru0_18; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1873 = _T_14 ? _GEN_1038 : plru0_19; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1874 = _T_14 ? _GEN_1039 : plru0_20; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1875 = _T_14 ? _GEN_1040 : plru0_21; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1876 = _T_14 ? _GEN_1041 : plru0_22; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1877 = _T_14 ? _GEN_1042 : plru0_23; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1878 = _T_14 ? _GEN_1043 : plru0_24; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1879 = _T_14 ? _GEN_1044 : plru0_25; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1880 = _T_14 ? _GEN_1045 : plru0_26; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1881 = _T_14 ? _GEN_1046 : plru0_27; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1882 = _T_14 ? _GEN_1047 : plru0_28; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1883 = _T_14 ? _GEN_1048 : plru0_29; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1884 = _T_14 ? _GEN_1049 : plru0_30; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1885 = _T_14 ? _GEN_1050 : plru0_31; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1886 = _T_14 ? _GEN_1051 : plru0_32; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1887 = _T_14 ? _GEN_1052 : plru0_33; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1888 = _T_14 ? _GEN_1053 : plru0_34; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1889 = _T_14 ? _GEN_1054 : plru0_35; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1890 = _T_14 ? _GEN_1055 : plru0_36; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1891 = _T_14 ? _GEN_1056 : plru0_37; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1892 = _T_14 ? _GEN_1057 : plru0_38; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1893 = _T_14 ? _GEN_1058 : plru0_39; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1894 = _T_14 ? _GEN_1059 : plru0_40; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1895 = _T_14 ? _GEN_1060 : plru0_41; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1896 = _T_14 ? _GEN_1061 : plru0_42; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1897 = _T_14 ? _GEN_1062 : plru0_43; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1898 = _T_14 ? _GEN_1063 : plru0_44; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1899 = _T_14 ? _GEN_1064 : plru0_45; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1900 = _T_14 ? _GEN_1065 : plru0_46; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1901 = _T_14 ? _GEN_1066 : plru0_47; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1902 = _T_14 ? _GEN_1067 : plru0_48; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1903 = _T_14 ? _GEN_1068 : plru0_49; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1904 = _T_14 ? _GEN_1069 : plru0_50; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1905 = _T_14 ? _GEN_1070 : plru0_51; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1906 = _T_14 ? _GEN_1071 : plru0_52; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1907 = _T_14 ? _GEN_1072 : plru0_53; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1908 = _T_14 ? _GEN_1073 : plru0_54; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1909 = _T_14 ? _GEN_1074 : plru0_55; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1910 = _T_14 ? _GEN_1075 : plru0_56; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1911 = _T_14 ? _GEN_1076 : plru0_57; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1912 = _T_14 ? _GEN_1077 : plru0_58; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1913 = _T_14 ? _GEN_1078 : plru0_59; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1914 = _T_14 ? _GEN_1079 : plru0_60; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1915 = _T_14 ? _GEN_1080 : plru0_61; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1916 = _T_14 ? _GEN_1081 : plru0_62; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1917 = _T_14 ? _GEN_1082 : plru0_63; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1918 = _T_14 ? _GEN_1211 : plru1_0; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1919 = _T_14 ? _GEN_1212 : plru1_1; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1920 = _T_14 ? _GEN_1213 : plru1_2; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1921 = _T_14 ? _GEN_1214 : plru1_3; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1922 = _T_14 ? _GEN_1215 : plru1_4; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1923 = _T_14 ? _GEN_1216 : plru1_5; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1924 = _T_14 ? _GEN_1217 : plru1_6; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1925 = _T_14 ? _GEN_1218 : plru1_7; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1926 = _T_14 ? _GEN_1219 : plru1_8; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1927 = _T_14 ? _GEN_1220 : plru1_9; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1928 = _T_14 ? _GEN_1221 : plru1_10; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1929 = _T_14 ? _GEN_1222 : plru1_11; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1930 = _T_14 ? _GEN_1223 : plru1_12; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1931 = _T_14 ? _GEN_1224 : plru1_13; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1932 = _T_14 ? _GEN_1225 : plru1_14; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1933 = _T_14 ? _GEN_1226 : plru1_15; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1934 = _T_14 ? _GEN_1227 : plru1_16; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1935 = _T_14 ? _GEN_1228 : plru1_17; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1936 = _T_14 ? _GEN_1229 : plru1_18; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1937 = _T_14 ? _GEN_1230 : plru1_19; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1938 = _T_14 ? _GEN_1231 : plru1_20; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1939 = _T_14 ? _GEN_1232 : plru1_21; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1940 = _T_14 ? _GEN_1233 : plru1_22; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1941 = _T_14 ? _GEN_1234 : plru1_23; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1942 = _T_14 ? _GEN_1235 : plru1_24; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1943 = _T_14 ? _GEN_1236 : plru1_25; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1944 = _T_14 ? _GEN_1237 : plru1_26; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1945 = _T_14 ? _GEN_1238 : plru1_27; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1946 = _T_14 ? _GEN_1239 : plru1_28; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1947 = _T_14 ? _GEN_1240 : plru1_29; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1948 = _T_14 ? _GEN_1241 : plru1_30; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1949 = _T_14 ? _GEN_1242 : plru1_31; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1950 = _T_14 ? _GEN_1243 : plru1_32; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1951 = _T_14 ? _GEN_1244 : plru1_33; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1952 = _T_14 ? _GEN_1245 : plru1_34; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1953 = _T_14 ? _GEN_1246 : plru1_35; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1954 = _T_14 ? _GEN_1247 : plru1_36; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1955 = _T_14 ? _GEN_1248 : plru1_37; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1956 = _T_14 ? _GEN_1249 : plru1_38; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1957 = _T_14 ? _GEN_1250 : plru1_39; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1958 = _T_14 ? _GEN_1251 : plru1_40; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1959 = _T_14 ? _GEN_1252 : plru1_41; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1960 = _T_14 ? _GEN_1253 : plru1_42; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1961 = _T_14 ? _GEN_1254 : plru1_43; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1962 = _T_14 ? _GEN_1255 : plru1_44; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1963 = _T_14 ? _GEN_1256 : plru1_45; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1964 = _T_14 ? _GEN_1257 : plru1_46; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1965 = _T_14 ? _GEN_1258 : plru1_47; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1966 = _T_14 ? _GEN_1259 : plru1_48; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1967 = _T_14 ? _GEN_1260 : plru1_49; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1968 = _T_14 ? _GEN_1261 : plru1_50; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1969 = _T_14 ? _GEN_1262 : plru1_51; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1970 = _T_14 ? _GEN_1263 : plru1_52; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1971 = _T_14 ? _GEN_1264 : plru1_53; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1972 = _T_14 ? _GEN_1265 : plru1_54; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1973 = _T_14 ? _GEN_1266 : plru1_55; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1974 = _T_14 ? _GEN_1267 : plru1_56; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1975 = _T_14 ? _GEN_1268 : plru1_57; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1976 = _T_14 ? _GEN_1269 : plru1_58; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1977 = _T_14 ? _GEN_1270 : plru1_59; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1978 = _T_14 ? _GEN_1271 : plru1_60; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1979 = _T_14 ? _GEN_1272 : plru1_61; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1980 = _T_14 ? _GEN_1273 : plru1_62; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1981 = _T_14 ? _GEN_1274 : plru1_63; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1982 = _T_14 ? _GEN_1275 : plru2_0; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1983 = _T_14 ? _GEN_1276 : plru2_1; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1984 = _T_14 ? _GEN_1277 : plru2_2; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1985 = _T_14 ? _GEN_1278 : plru2_3; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1986 = _T_14 ? _GEN_1279 : plru2_4; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1987 = _T_14 ? _GEN_1280 : plru2_5; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1988 = _T_14 ? _GEN_1281 : plru2_6; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1989 = _T_14 ? _GEN_1282 : plru2_7; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1990 = _T_14 ? _GEN_1283 : plru2_8; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1991 = _T_14 ? _GEN_1284 : plru2_9; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1992 = _T_14 ? _GEN_1285 : plru2_10; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1993 = _T_14 ? _GEN_1286 : plru2_11; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1994 = _T_14 ? _GEN_1287 : plru2_12; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1995 = _T_14 ? _GEN_1288 : plru2_13; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1996 = _T_14 ? _GEN_1289 : plru2_14; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1997 = _T_14 ? _GEN_1290 : plru2_15; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1998 = _T_14 ? _GEN_1291 : plru2_16; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1999 = _T_14 ? _GEN_1292 : plru2_17; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2000 = _T_14 ? _GEN_1293 : plru2_18; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2001 = _T_14 ? _GEN_1294 : plru2_19; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2002 = _T_14 ? _GEN_1295 : plru2_20; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2003 = _T_14 ? _GEN_1296 : plru2_21; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2004 = _T_14 ? _GEN_1297 : plru2_22; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2005 = _T_14 ? _GEN_1298 : plru2_23; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2006 = _T_14 ? _GEN_1299 : plru2_24; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2007 = _T_14 ? _GEN_1300 : plru2_25; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2008 = _T_14 ? _GEN_1301 : plru2_26; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2009 = _T_14 ? _GEN_1302 : plru2_27; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2010 = _T_14 ? _GEN_1303 : plru2_28; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2011 = _T_14 ? _GEN_1304 : plru2_29; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2012 = _T_14 ? _GEN_1305 : plru2_30; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2013 = _T_14 ? _GEN_1306 : plru2_31; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2014 = _T_14 ? _GEN_1307 : plru2_32; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2015 = _T_14 ? _GEN_1308 : plru2_33; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2016 = _T_14 ? _GEN_1309 : plru2_34; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2017 = _T_14 ? _GEN_1310 : plru2_35; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2018 = _T_14 ? _GEN_1311 : plru2_36; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2019 = _T_14 ? _GEN_1312 : plru2_37; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2020 = _T_14 ? _GEN_1313 : plru2_38; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2021 = _T_14 ? _GEN_1314 : plru2_39; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2022 = _T_14 ? _GEN_1315 : plru2_40; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2023 = _T_14 ? _GEN_1316 : plru2_41; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2024 = _T_14 ? _GEN_1317 : plru2_42; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2025 = _T_14 ? _GEN_1318 : plru2_43; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2026 = _T_14 ? _GEN_1319 : plru2_44; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2027 = _T_14 ? _GEN_1320 : plru2_45; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2028 = _T_14 ? _GEN_1321 : plru2_46; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2029 = _T_14 ? _GEN_1322 : plru2_47; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2030 = _T_14 ? _GEN_1323 : plru2_48; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2031 = _T_14 ? _GEN_1324 : plru2_49; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2032 = _T_14 ? _GEN_1325 : plru2_50; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2033 = _T_14 ? _GEN_1326 : plru2_51; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2034 = _T_14 ? _GEN_1327 : plru2_52; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2035 = _T_14 ? _GEN_1328 : plru2_53; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2036 = _T_14 ? _GEN_1329 : plru2_54; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2037 = _T_14 ? _GEN_1330 : plru2_55; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2038 = _T_14 ? _GEN_1331 : plru2_56; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2039 = _T_14 ? _GEN_1332 : plru2_57; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2040 = _T_14 ? _GEN_1333 : plru2_58; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2041 = _T_14 ? _GEN_1334 : plru2_59; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2042 = _T_14 ? _GEN_1335 : plru2_60; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2043 = _T_14 ? _GEN_1336 : plru2_61; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2044 = _T_14 ? _GEN_1337 : plru2_62; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2045 = _T_14 ? _GEN_1338 : plru2_63; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire [3:0] _GEN_2046 = _T_14 ? 4'h7 : state; // @[Cache.scala 368:30 Cache.scala 370:15 Cache.scala 207:22]
  wire  _T_31 = 4'h7 == state; // @[Conditional.scala 37:30]
  reg [63:0] io_in_resp_bits_rdata_REG; // @[Cache.scala 374:36]
  wire  _T_32 = io_in_resp_ready & io_in_resp_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_2047 = _T_32 ? 4'h8 : state; // @[Cache.scala 375:29 Cache.scala 376:15 Cache.scala 207:22]
  wire [63:0] _GEN_2048 = _T_31 ? io_in_resp_bits_rdata_REG : 64'h0; // @[Conditional.scala 39:67 Cache.scala 374:26 Cache.scala 277:22]
  wire [3:0] _GEN_2049 = _T_31 ? _GEN_2047 : state; // @[Conditional.scala 39:67 Cache.scala 207:22]
  wire  _GEN_2050 = _T_27 ? 1'h0 : _GEN_27; // @[Conditional.scala 39:67 Cache.scala 367:14]
  wire  _GEN_2051 = _T_27 ? _GEN_1854 : plru0_0; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2052 = _T_27 ? _GEN_1855 : plru0_1; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2053 = _T_27 ? _GEN_1856 : plru0_2; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2054 = _T_27 ? _GEN_1857 : plru0_3; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2055 = _T_27 ? _GEN_1858 : plru0_4; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2056 = _T_27 ? _GEN_1859 : plru0_5; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2057 = _T_27 ? _GEN_1860 : plru0_6; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2058 = _T_27 ? _GEN_1861 : plru0_7; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2059 = _T_27 ? _GEN_1862 : plru0_8; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2060 = _T_27 ? _GEN_1863 : plru0_9; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2061 = _T_27 ? _GEN_1864 : plru0_10; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2062 = _T_27 ? _GEN_1865 : plru0_11; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2063 = _T_27 ? _GEN_1866 : plru0_12; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2064 = _T_27 ? _GEN_1867 : plru0_13; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2065 = _T_27 ? _GEN_1868 : plru0_14; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2066 = _T_27 ? _GEN_1869 : plru0_15; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2067 = _T_27 ? _GEN_1870 : plru0_16; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2068 = _T_27 ? _GEN_1871 : plru0_17; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2069 = _T_27 ? _GEN_1872 : plru0_18; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2070 = _T_27 ? _GEN_1873 : plru0_19; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2071 = _T_27 ? _GEN_1874 : plru0_20; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2072 = _T_27 ? _GEN_1875 : plru0_21; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2073 = _T_27 ? _GEN_1876 : plru0_22; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2074 = _T_27 ? _GEN_1877 : plru0_23; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2075 = _T_27 ? _GEN_1878 : plru0_24; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2076 = _T_27 ? _GEN_1879 : plru0_25; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2077 = _T_27 ? _GEN_1880 : plru0_26; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2078 = _T_27 ? _GEN_1881 : plru0_27; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2079 = _T_27 ? _GEN_1882 : plru0_28; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2080 = _T_27 ? _GEN_1883 : plru0_29; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2081 = _T_27 ? _GEN_1884 : plru0_30; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2082 = _T_27 ? _GEN_1885 : plru0_31; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2083 = _T_27 ? _GEN_1886 : plru0_32; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2084 = _T_27 ? _GEN_1887 : plru0_33; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2085 = _T_27 ? _GEN_1888 : plru0_34; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2086 = _T_27 ? _GEN_1889 : plru0_35; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2087 = _T_27 ? _GEN_1890 : plru0_36; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2088 = _T_27 ? _GEN_1891 : plru0_37; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2089 = _T_27 ? _GEN_1892 : plru0_38; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2090 = _T_27 ? _GEN_1893 : plru0_39; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2091 = _T_27 ? _GEN_1894 : plru0_40; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2092 = _T_27 ? _GEN_1895 : plru0_41; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2093 = _T_27 ? _GEN_1896 : plru0_42; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2094 = _T_27 ? _GEN_1897 : plru0_43; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2095 = _T_27 ? _GEN_1898 : plru0_44; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2096 = _T_27 ? _GEN_1899 : plru0_45; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2097 = _T_27 ? _GEN_1900 : plru0_46; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2098 = _T_27 ? _GEN_1901 : plru0_47; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2099 = _T_27 ? _GEN_1902 : plru0_48; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2100 = _T_27 ? _GEN_1903 : plru0_49; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2101 = _T_27 ? _GEN_1904 : plru0_50; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2102 = _T_27 ? _GEN_1905 : plru0_51; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2103 = _T_27 ? _GEN_1906 : plru0_52; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2104 = _T_27 ? _GEN_1907 : plru0_53; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2105 = _T_27 ? _GEN_1908 : plru0_54; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2106 = _T_27 ? _GEN_1909 : plru0_55; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2107 = _T_27 ? _GEN_1910 : plru0_56; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2108 = _T_27 ? _GEN_1911 : plru0_57; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2109 = _T_27 ? _GEN_1912 : plru0_58; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2110 = _T_27 ? _GEN_1913 : plru0_59; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2111 = _T_27 ? _GEN_1914 : plru0_60; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2112 = _T_27 ? _GEN_1915 : plru0_61; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2113 = _T_27 ? _GEN_1916 : plru0_62; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2114 = _T_27 ? _GEN_1917 : plru0_63; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2115 = _T_27 ? _GEN_1918 : plru1_0; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2116 = _T_27 ? _GEN_1919 : plru1_1; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2117 = _T_27 ? _GEN_1920 : plru1_2; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2118 = _T_27 ? _GEN_1921 : plru1_3; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2119 = _T_27 ? _GEN_1922 : plru1_4; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2120 = _T_27 ? _GEN_1923 : plru1_5; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2121 = _T_27 ? _GEN_1924 : plru1_6; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2122 = _T_27 ? _GEN_1925 : plru1_7; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2123 = _T_27 ? _GEN_1926 : plru1_8; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2124 = _T_27 ? _GEN_1927 : plru1_9; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2125 = _T_27 ? _GEN_1928 : plru1_10; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2126 = _T_27 ? _GEN_1929 : plru1_11; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2127 = _T_27 ? _GEN_1930 : plru1_12; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2128 = _T_27 ? _GEN_1931 : plru1_13; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2129 = _T_27 ? _GEN_1932 : plru1_14; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2130 = _T_27 ? _GEN_1933 : plru1_15; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2131 = _T_27 ? _GEN_1934 : plru1_16; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2132 = _T_27 ? _GEN_1935 : plru1_17; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2133 = _T_27 ? _GEN_1936 : plru1_18; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2134 = _T_27 ? _GEN_1937 : plru1_19; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2135 = _T_27 ? _GEN_1938 : plru1_20; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2136 = _T_27 ? _GEN_1939 : plru1_21; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2137 = _T_27 ? _GEN_1940 : plru1_22; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2138 = _T_27 ? _GEN_1941 : plru1_23; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2139 = _T_27 ? _GEN_1942 : plru1_24; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2140 = _T_27 ? _GEN_1943 : plru1_25; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2141 = _T_27 ? _GEN_1944 : plru1_26; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2142 = _T_27 ? _GEN_1945 : plru1_27; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2143 = _T_27 ? _GEN_1946 : plru1_28; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2144 = _T_27 ? _GEN_1947 : plru1_29; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2145 = _T_27 ? _GEN_1948 : plru1_30; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2146 = _T_27 ? _GEN_1949 : plru1_31; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2147 = _T_27 ? _GEN_1950 : plru1_32; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2148 = _T_27 ? _GEN_1951 : plru1_33; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2149 = _T_27 ? _GEN_1952 : plru1_34; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2150 = _T_27 ? _GEN_1953 : plru1_35; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2151 = _T_27 ? _GEN_1954 : plru1_36; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2152 = _T_27 ? _GEN_1955 : plru1_37; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2153 = _T_27 ? _GEN_1956 : plru1_38; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2154 = _T_27 ? _GEN_1957 : plru1_39; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2155 = _T_27 ? _GEN_1958 : plru1_40; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2156 = _T_27 ? _GEN_1959 : plru1_41; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2157 = _T_27 ? _GEN_1960 : plru1_42; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2158 = _T_27 ? _GEN_1961 : plru1_43; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2159 = _T_27 ? _GEN_1962 : plru1_44; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2160 = _T_27 ? _GEN_1963 : plru1_45; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2161 = _T_27 ? _GEN_1964 : plru1_46; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2162 = _T_27 ? _GEN_1965 : plru1_47; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2163 = _T_27 ? _GEN_1966 : plru1_48; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2164 = _T_27 ? _GEN_1967 : plru1_49; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2165 = _T_27 ? _GEN_1968 : plru1_50; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2166 = _T_27 ? _GEN_1969 : plru1_51; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2167 = _T_27 ? _GEN_1970 : plru1_52; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2168 = _T_27 ? _GEN_1971 : plru1_53; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2169 = _T_27 ? _GEN_1972 : plru1_54; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2170 = _T_27 ? _GEN_1973 : plru1_55; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2171 = _T_27 ? _GEN_1974 : plru1_56; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2172 = _T_27 ? _GEN_1975 : plru1_57; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2173 = _T_27 ? _GEN_1976 : plru1_58; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2174 = _T_27 ? _GEN_1977 : plru1_59; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2175 = _T_27 ? _GEN_1978 : plru1_60; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2176 = _T_27 ? _GEN_1979 : plru1_61; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2177 = _T_27 ? _GEN_1980 : plru1_62; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2178 = _T_27 ? _GEN_1981 : plru1_63; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2179 = _T_27 ? _GEN_1982 : plru2_0; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2180 = _T_27 ? _GEN_1983 : plru2_1; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2181 = _T_27 ? _GEN_1984 : plru2_2; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2182 = _T_27 ? _GEN_1985 : plru2_3; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2183 = _T_27 ? _GEN_1986 : plru2_4; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2184 = _T_27 ? _GEN_1987 : plru2_5; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2185 = _T_27 ? _GEN_1988 : plru2_6; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2186 = _T_27 ? _GEN_1989 : plru2_7; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2187 = _T_27 ? _GEN_1990 : plru2_8; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2188 = _T_27 ? _GEN_1991 : plru2_9; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2189 = _T_27 ? _GEN_1992 : plru2_10; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2190 = _T_27 ? _GEN_1993 : plru2_11; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2191 = _T_27 ? _GEN_1994 : plru2_12; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2192 = _T_27 ? _GEN_1995 : plru2_13; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2193 = _T_27 ? _GEN_1996 : plru2_14; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2194 = _T_27 ? _GEN_1997 : plru2_15; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2195 = _T_27 ? _GEN_1998 : plru2_16; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2196 = _T_27 ? _GEN_1999 : plru2_17; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2197 = _T_27 ? _GEN_2000 : plru2_18; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2198 = _T_27 ? _GEN_2001 : plru2_19; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2199 = _T_27 ? _GEN_2002 : plru2_20; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2200 = _T_27 ? _GEN_2003 : plru2_21; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2201 = _T_27 ? _GEN_2004 : plru2_22; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2202 = _T_27 ? _GEN_2005 : plru2_23; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2203 = _T_27 ? _GEN_2006 : plru2_24; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2204 = _T_27 ? _GEN_2007 : plru2_25; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2205 = _T_27 ? _GEN_2008 : plru2_26; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2206 = _T_27 ? _GEN_2009 : plru2_27; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2207 = _T_27 ? _GEN_2010 : plru2_28; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2208 = _T_27 ? _GEN_2011 : plru2_29; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2209 = _T_27 ? _GEN_2012 : plru2_30; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2210 = _T_27 ? _GEN_2013 : plru2_31; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2211 = _T_27 ? _GEN_2014 : plru2_32; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2212 = _T_27 ? _GEN_2015 : plru2_33; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2213 = _T_27 ? _GEN_2016 : plru2_34; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2214 = _T_27 ? _GEN_2017 : plru2_35; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2215 = _T_27 ? _GEN_2018 : plru2_36; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2216 = _T_27 ? _GEN_2019 : plru2_37; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2217 = _T_27 ? _GEN_2020 : plru2_38; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2218 = _T_27 ? _GEN_2021 : plru2_39; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2219 = _T_27 ? _GEN_2022 : plru2_40; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2220 = _T_27 ? _GEN_2023 : plru2_41; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2221 = _T_27 ? _GEN_2024 : plru2_42; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2222 = _T_27 ? _GEN_2025 : plru2_43; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2223 = _T_27 ? _GEN_2026 : plru2_44; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2224 = _T_27 ? _GEN_2027 : plru2_45; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2225 = _T_27 ? _GEN_2028 : plru2_46; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2226 = _T_27 ? _GEN_2029 : plru2_47; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2227 = _T_27 ? _GEN_2030 : plru2_48; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2228 = _T_27 ? _GEN_2031 : plru2_49; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2229 = _T_27 ? _GEN_2032 : plru2_50; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2230 = _T_27 ? _GEN_2033 : plru2_51; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2231 = _T_27 ? _GEN_2034 : plru2_52; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2232 = _T_27 ? _GEN_2035 : plru2_53; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2233 = _T_27 ? _GEN_2036 : plru2_54; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2234 = _T_27 ? _GEN_2037 : plru2_55; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2235 = _T_27 ? _GEN_2038 : plru2_56; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2236 = _T_27 ? _GEN_2039 : plru2_57; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2237 = _T_27 ? _GEN_2040 : plru2_58; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2238 = _T_27 ? _GEN_2041 : plru2_59; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2239 = _T_27 ? _GEN_2042 : plru2_60; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2240 = _T_27 ? _GEN_2043 : plru2_61; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2241 = _T_27 ? _GEN_2044 : plru2_62; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2242 = _T_27 ? _GEN_2045 : plru2_63; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire [3:0] _GEN_2243 = _T_27 ? _GEN_2046 : _GEN_2049; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_2244 = _T_27 ? 64'h0 : _GEN_2048; // @[Conditional.scala 39:67 Cache.scala 277:22]
  wire [3:0] _GEN_2245 = _T_25 ? _GEN_1533 : _GEN_2243; // @[Conditional.scala 39:67]
  wire  _GEN_2246 = _T_25 ? _GEN_27 : _GEN_2050; // @[Conditional.scala 39:67]
  wire  _GEN_2247 = _T_25 ? plru0_0 : _GEN_2051; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2248 = _T_25 ? plru0_1 : _GEN_2052; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2249 = _T_25 ? plru0_2 : _GEN_2053; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2250 = _T_25 ? plru0_3 : _GEN_2054; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2251 = _T_25 ? plru0_4 : _GEN_2055; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2252 = _T_25 ? plru0_5 : _GEN_2056; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2253 = _T_25 ? plru0_6 : _GEN_2057; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2254 = _T_25 ? plru0_7 : _GEN_2058; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2255 = _T_25 ? plru0_8 : _GEN_2059; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2256 = _T_25 ? plru0_9 : _GEN_2060; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2257 = _T_25 ? plru0_10 : _GEN_2061; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2258 = _T_25 ? plru0_11 : _GEN_2062; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2259 = _T_25 ? plru0_12 : _GEN_2063; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2260 = _T_25 ? plru0_13 : _GEN_2064; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2261 = _T_25 ? plru0_14 : _GEN_2065; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2262 = _T_25 ? plru0_15 : _GEN_2066; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2263 = _T_25 ? plru0_16 : _GEN_2067; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2264 = _T_25 ? plru0_17 : _GEN_2068; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2265 = _T_25 ? plru0_18 : _GEN_2069; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2266 = _T_25 ? plru0_19 : _GEN_2070; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2267 = _T_25 ? plru0_20 : _GEN_2071; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2268 = _T_25 ? plru0_21 : _GEN_2072; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2269 = _T_25 ? plru0_22 : _GEN_2073; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2270 = _T_25 ? plru0_23 : _GEN_2074; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2271 = _T_25 ? plru0_24 : _GEN_2075; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2272 = _T_25 ? plru0_25 : _GEN_2076; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2273 = _T_25 ? plru0_26 : _GEN_2077; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2274 = _T_25 ? plru0_27 : _GEN_2078; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2275 = _T_25 ? plru0_28 : _GEN_2079; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2276 = _T_25 ? plru0_29 : _GEN_2080; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2277 = _T_25 ? plru0_30 : _GEN_2081; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2278 = _T_25 ? plru0_31 : _GEN_2082; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2279 = _T_25 ? plru0_32 : _GEN_2083; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2280 = _T_25 ? plru0_33 : _GEN_2084; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2281 = _T_25 ? plru0_34 : _GEN_2085; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2282 = _T_25 ? plru0_35 : _GEN_2086; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2283 = _T_25 ? plru0_36 : _GEN_2087; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2284 = _T_25 ? plru0_37 : _GEN_2088; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2285 = _T_25 ? plru0_38 : _GEN_2089; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2286 = _T_25 ? plru0_39 : _GEN_2090; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2287 = _T_25 ? plru0_40 : _GEN_2091; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2288 = _T_25 ? plru0_41 : _GEN_2092; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2289 = _T_25 ? plru0_42 : _GEN_2093; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2290 = _T_25 ? plru0_43 : _GEN_2094; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2291 = _T_25 ? plru0_44 : _GEN_2095; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2292 = _T_25 ? plru0_45 : _GEN_2096; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2293 = _T_25 ? plru0_46 : _GEN_2097; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2294 = _T_25 ? plru0_47 : _GEN_2098; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2295 = _T_25 ? plru0_48 : _GEN_2099; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2296 = _T_25 ? plru0_49 : _GEN_2100; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2297 = _T_25 ? plru0_50 : _GEN_2101; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2298 = _T_25 ? plru0_51 : _GEN_2102; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2299 = _T_25 ? plru0_52 : _GEN_2103; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2300 = _T_25 ? plru0_53 : _GEN_2104; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2301 = _T_25 ? plru0_54 : _GEN_2105; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2302 = _T_25 ? plru0_55 : _GEN_2106; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2303 = _T_25 ? plru0_56 : _GEN_2107; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2304 = _T_25 ? plru0_57 : _GEN_2108; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2305 = _T_25 ? plru0_58 : _GEN_2109; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2306 = _T_25 ? plru0_59 : _GEN_2110; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2307 = _T_25 ? plru0_60 : _GEN_2111; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2308 = _T_25 ? plru0_61 : _GEN_2112; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2309 = _T_25 ? plru0_62 : _GEN_2113; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2310 = _T_25 ? plru0_63 : _GEN_2114; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2311 = _T_25 ? plru1_0 : _GEN_2115; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2312 = _T_25 ? plru1_1 : _GEN_2116; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2313 = _T_25 ? plru1_2 : _GEN_2117; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2314 = _T_25 ? plru1_3 : _GEN_2118; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2315 = _T_25 ? plru1_4 : _GEN_2119; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2316 = _T_25 ? plru1_5 : _GEN_2120; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2317 = _T_25 ? plru1_6 : _GEN_2121; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2318 = _T_25 ? plru1_7 : _GEN_2122; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2319 = _T_25 ? plru1_8 : _GEN_2123; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2320 = _T_25 ? plru1_9 : _GEN_2124; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2321 = _T_25 ? plru1_10 : _GEN_2125; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2322 = _T_25 ? plru1_11 : _GEN_2126; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2323 = _T_25 ? plru1_12 : _GEN_2127; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2324 = _T_25 ? plru1_13 : _GEN_2128; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2325 = _T_25 ? plru1_14 : _GEN_2129; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2326 = _T_25 ? plru1_15 : _GEN_2130; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2327 = _T_25 ? plru1_16 : _GEN_2131; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2328 = _T_25 ? plru1_17 : _GEN_2132; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2329 = _T_25 ? plru1_18 : _GEN_2133; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2330 = _T_25 ? plru1_19 : _GEN_2134; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2331 = _T_25 ? plru1_20 : _GEN_2135; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2332 = _T_25 ? plru1_21 : _GEN_2136; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2333 = _T_25 ? plru1_22 : _GEN_2137; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2334 = _T_25 ? plru1_23 : _GEN_2138; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2335 = _T_25 ? plru1_24 : _GEN_2139; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2336 = _T_25 ? plru1_25 : _GEN_2140; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2337 = _T_25 ? plru1_26 : _GEN_2141; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2338 = _T_25 ? plru1_27 : _GEN_2142; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2339 = _T_25 ? plru1_28 : _GEN_2143; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2340 = _T_25 ? plru1_29 : _GEN_2144; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2341 = _T_25 ? plru1_30 : _GEN_2145; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2342 = _T_25 ? plru1_31 : _GEN_2146; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2343 = _T_25 ? plru1_32 : _GEN_2147; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2344 = _T_25 ? plru1_33 : _GEN_2148; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2345 = _T_25 ? plru1_34 : _GEN_2149; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2346 = _T_25 ? plru1_35 : _GEN_2150; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2347 = _T_25 ? plru1_36 : _GEN_2151; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2348 = _T_25 ? plru1_37 : _GEN_2152; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2349 = _T_25 ? plru1_38 : _GEN_2153; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2350 = _T_25 ? plru1_39 : _GEN_2154; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2351 = _T_25 ? plru1_40 : _GEN_2155; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2352 = _T_25 ? plru1_41 : _GEN_2156; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2353 = _T_25 ? plru1_42 : _GEN_2157; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2354 = _T_25 ? plru1_43 : _GEN_2158; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2355 = _T_25 ? plru1_44 : _GEN_2159; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2356 = _T_25 ? plru1_45 : _GEN_2160; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2357 = _T_25 ? plru1_46 : _GEN_2161; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2358 = _T_25 ? plru1_47 : _GEN_2162; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2359 = _T_25 ? plru1_48 : _GEN_2163; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2360 = _T_25 ? plru1_49 : _GEN_2164; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2361 = _T_25 ? plru1_50 : _GEN_2165; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2362 = _T_25 ? plru1_51 : _GEN_2166; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2363 = _T_25 ? plru1_52 : _GEN_2167; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2364 = _T_25 ? plru1_53 : _GEN_2168; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2365 = _T_25 ? plru1_54 : _GEN_2169; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2366 = _T_25 ? plru1_55 : _GEN_2170; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2367 = _T_25 ? plru1_56 : _GEN_2171; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2368 = _T_25 ? plru1_57 : _GEN_2172; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2369 = _T_25 ? plru1_58 : _GEN_2173; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2370 = _T_25 ? plru1_59 : _GEN_2174; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2371 = _T_25 ? plru1_60 : _GEN_2175; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2372 = _T_25 ? plru1_61 : _GEN_2176; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2373 = _T_25 ? plru1_62 : _GEN_2177; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2374 = _T_25 ? plru1_63 : _GEN_2178; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2375 = _T_25 ? plru2_0 : _GEN_2179; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2376 = _T_25 ? plru2_1 : _GEN_2180; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2377 = _T_25 ? plru2_2 : _GEN_2181; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2378 = _T_25 ? plru2_3 : _GEN_2182; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2379 = _T_25 ? plru2_4 : _GEN_2183; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2380 = _T_25 ? plru2_5 : _GEN_2184; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2381 = _T_25 ? plru2_6 : _GEN_2185; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2382 = _T_25 ? plru2_7 : _GEN_2186; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2383 = _T_25 ? plru2_8 : _GEN_2187; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2384 = _T_25 ? plru2_9 : _GEN_2188; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2385 = _T_25 ? plru2_10 : _GEN_2189; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2386 = _T_25 ? plru2_11 : _GEN_2190; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2387 = _T_25 ? plru2_12 : _GEN_2191; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2388 = _T_25 ? plru2_13 : _GEN_2192; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2389 = _T_25 ? plru2_14 : _GEN_2193; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2390 = _T_25 ? plru2_15 : _GEN_2194; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2391 = _T_25 ? plru2_16 : _GEN_2195; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2392 = _T_25 ? plru2_17 : _GEN_2196; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2393 = _T_25 ? plru2_18 : _GEN_2197; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2394 = _T_25 ? plru2_19 : _GEN_2198; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2395 = _T_25 ? plru2_20 : _GEN_2199; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2396 = _T_25 ? plru2_21 : _GEN_2200; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2397 = _T_25 ? plru2_22 : _GEN_2201; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2398 = _T_25 ? plru2_23 : _GEN_2202; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2399 = _T_25 ? plru2_24 : _GEN_2203; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2400 = _T_25 ? plru2_25 : _GEN_2204; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2401 = _T_25 ? plru2_26 : _GEN_2205; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2402 = _T_25 ? plru2_27 : _GEN_2206; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2403 = _T_25 ? plru2_28 : _GEN_2207; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2404 = _T_25 ? plru2_29 : _GEN_2208; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2405 = _T_25 ? plru2_30 : _GEN_2209; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2406 = _T_25 ? plru2_31 : _GEN_2210; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2407 = _T_25 ? plru2_32 : _GEN_2211; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2408 = _T_25 ? plru2_33 : _GEN_2212; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2409 = _T_25 ? plru2_34 : _GEN_2213; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2410 = _T_25 ? plru2_35 : _GEN_2214; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2411 = _T_25 ? plru2_36 : _GEN_2215; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2412 = _T_25 ? plru2_37 : _GEN_2216; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2413 = _T_25 ? plru2_38 : _GEN_2217; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2414 = _T_25 ? plru2_39 : _GEN_2218; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2415 = _T_25 ? plru2_40 : _GEN_2219; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2416 = _T_25 ? plru2_41 : _GEN_2220; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2417 = _T_25 ? plru2_42 : _GEN_2221; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2418 = _T_25 ? plru2_43 : _GEN_2222; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2419 = _T_25 ? plru2_44 : _GEN_2223; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2420 = _T_25 ? plru2_45 : _GEN_2224; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2421 = _T_25 ? plru2_46 : _GEN_2225; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2422 = _T_25 ? plru2_47 : _GEN_2226; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2423 = _T_25 ? plru2_48 : _GEN_2227; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2424 = _T_25 ? plru2_49 : _GEN_2228; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2425 = _T_25 ? plru2_50 : _GEN_2229; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2426 = _T_25 ? plru2_51 : _GEN_2230; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2427 = _T_25 ? plru2_52 : _GEN_2231; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2428 = _T_25 ? plru2_53 : _GEN_2232; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2429 = _T_25 ? plru2_54 : _GEN_2233; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2430 = _T_25 ? plru2_55 : _GEN_2234; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2431 = _T_25 ? plru2_56 : _GEN_2235; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2432 = _T_25 ? plru2_57 : _GEN_2236; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2433 = _T_25 ? plru2_58 : _GEN_2237; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2434 = _T_25 ? plru2_59 : _GEN_2238; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2435 = _T_25 ? plru2_60 : _GEN_2239; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2436 = _T_25 ? plru2_61 : _GEN_2240; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2437 = _T_25 ? plru2_62 : _GEN_2241; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2438 = _T_25 ? plru2_63 : _GEN_2242; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire [63:0] _GEN_2439 = _T_25 ? 64'h0 : _GEN_2244; // @[Conditional.scala 39:67 Cache.scala 277:22]
  wire [3:0] _GEN_2440 = _T_23 ? _GEN_1532 : _GEN_2245; // @[Conditional.scala 39:67]
  wire  _GEN_2441 = _T_23 ? _GEN_27 : _GEN_2246; // @[Conditional.scala 39:67]
  wire  _GEN_2442 = _T_23 ? plru0_0 : _GEN_2247; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2443 = _T_23 ? plru0_1 : _GEN_2248; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2444 = _T_23 ? plru0_2 : _GEN_2249; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2445 = _T_23 ? plru0_3 : _GEN_2250; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2446 = _T_23 ? plru0_4 : _GEN_2251; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2447 = _T_23 ? plru0_5 : _GEN_2252; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2448 = _T_23 ? plru0_6 : _GEN_2253; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2449 = _T_23 ? plru0_7 : _GEN_2254; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2450 = _T_23 ? plru0_8 : _GEN_2255; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2451 = _T_23 ? plru0_9 : _GEN_2256; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2452 = _T_23 ? plru0_10 : _GEN_2257; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2453 = _T_23 ? plru0_11 : _GEN_2258; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2454 = _T_23 ? plru0_12 : _GEN_2259; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2455 = _T_23 ? plru0_13 : _GEN_2260; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2456 = _T_23 ? plru0_14 : _GEN_2261; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2457 = _T_23 ? plru0_15 : _GEN_2262; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2458 = _T_23 ? plru0_16 : _GEN_2263; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2459 = _T_23 ? plru0_17 : _GEN_2264; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2460 = _T_23 ? plru0_18 : _GEN_2265; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2461 = _T_23 ? plru0_19 : _GEN_2266; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2462 = _T_23 ? plru0_20 : _GEN_2267; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2463 = _T_23 ? plru0_21 : _GEN_2268; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2464 = _T_23 ? plru0_22 : _GEN_2269; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2465 = _T_23 ? plru0_23 : _GEN_2270; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2466 = _T_23 ? plru0_24 : _GEN_2271; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2467 = _T_23 ? plru0_25 : _GEN_2272; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2468 = _T_23 ? plru0_26 : _GEN_2273; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2469 = _T_23 ? plru0_27 : _GEN_2274; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2470 = _T_23 ? plru0_28 : _GEN_2275; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2471 = _T_23 ? plru0_29 : _GEN_2276; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2472 = _T_23 ? plru0_30 : _GEN_2277; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2473 = _T_23 ? plru0_31 : _GEN_2278; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2474 = _T_23 ? plru0_32 : _GEN_2279; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2475 = _T_23 ? plru0_33 : _GEN_2280; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2476 = _T_23 ? plru0_34 : _GEN_2281; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2477 = _T_23 ? plru0_35 : _GEN_2282; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2478 = _T_23 ? plru0_36 : _GEN_2283; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2479 = _T_23 ? plru0_37 : _GEN_2284; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2480 = _T_23 ? plru0_38 : _GEN_2285; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2481 = _T_23 ? plru0_39 : _GEN_2286; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2482 = _T_23 ? plru0_40 : _GEN_2287; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2483 = _T_23 ? plru0_41 : _GEN_2288; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2484 = _T_23 ? plru0_42 : _GEN_2289; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2485 = _T_23 ? plru0_43 : _GEN_2290; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2486 = _T_23 ? plru0_44 : _GEN_2291; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2487 = _T_23 ? plru0_45 : _GEN_2292; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2488 = _T_23 ? plru0_46 : _GEN_2293; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2489 = _T_23 ? plru0_47 : _GEN_2294; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2490 = _T_23 ? plru0_48 : _GEN_2295; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2491 = _T_23 ? plru0_49 : _GEN_2296; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2492 = _T_23 ? plru0_50 : _GEN_2297; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2493 = _T_23 ? plru0_51 : _GEN_2298; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2494 = _T_23 ? plru0_52 : _GEN_2299; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2495 = _T_23 ? plru0_53 : _GEN_2300; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2496 = _T_23 ? plru0_54 : _GEN_2301; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2497 = _T_23 ? plru0_55 : _GEN_2302; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2498 = _T_23 ? plru0_56 : _GEN_2303; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2499 = _T_23 ? plru0_57 : _GEN_2304; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2500 = _T_23 ? plru0_58 : _GEN_2305; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2501 = _T_23 ? plru0_59 : _GEN_2306; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2502 = _T_23 ? plru0_60 : _GEN_2307; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2503 = _T_23 ? plru0_61 : _GEN_2308; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2504 = _T_23 ? plru0_62 : _GEN_2309; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2505 = _T_23 ? plru0_63 : _GEN_2310; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2506 = _T_23 ? plru1_0 : _GEN_2311; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2507 = _T_23 ? plru1_1 : _GEN_2312; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2508 = _T_23 ? plru1_2 : _GEN_2313; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2509 = _T_23 ? plru1_3 : _GEN_2314; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2510 = _T_23 ? plru1_4 : _GEN_2315; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2511 = _T_23 ? plru1_5 : _GEN_2316; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2512 = _T_23 ? plru1_6 : _GEN_2317; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2513 = _T_23 ? plru1_7 : _GEN_2318; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2514 = _T_23 ? plru1_8 : _GEN_2319; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2515 = _T_23 ? plru1_9 : _GEN_2320; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2516 = _T_23 ? plru1_10 : _GEN_2321; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2517 = _T_23 ? plru1_11 : _GEN_2322; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2518 = _T_23 ? plru1_12 : _GEN_2323; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2519 = _T_23 ? plru1_13 : _GEN_2324; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2520 = _T_23 ? plru1_14 : _GEN_2325; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2521 = _T_23 ? plru1_15 : _GEN_2326; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2522 = _T_23 ? plru1_16 : _GEN_2327; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2523 = _T_23 ? plru1_17 : _GEN_2328; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2524 = _T_23 ? plru1_18 : _GEN_2329; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2525 = _T_23 ? plru1_19 : _GEN_2330; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2526 = _T_23 ? plru1_20 : _GEN_2331; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2527 = _T_23 ? plru1_21 : _GEN_2332; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2528 = _T_23 ? plru1_22 : _GEN_2333; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2529 = _T_23 ? plru1_23 : _GEN_2334; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2530 = _T_23 ? plru1_24 : _GEN_2335; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2531 = _T_23 ? plru1_25 : _GEN_2336; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2532 = _T_23 ? plru1_26 : _GEN_2337; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2533 = _T_23 ? plru1_27 : _GEN_2338; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2534 = _T_23 ? plru1_28 : _GEN_2339; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2535 = _T_23 ? plru1_29 : _GEN_2340; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2536 = _T_23 ? plru1_30 : _GEN_2341; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2537 = _T_23 ? plru1_31 : _GEN_2342; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2538 = _T_23 ? plru1_32 : _GEN_2343; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2539 = _T_23 ? plru1_33 : _GEN_2344; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2540 = _T_23 ? plru1_34 : _GEN_2345; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2541 = _T_23 ? plru1_35 : _GEN_2346; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2542 = _T_23 ? plru1_36 : _GEN_2347; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2543 = _T_23 ? plru1_37 : _GEN_2348; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2544 = _T_23 ? plru1_38 : _GEN_2349; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2545 = _T_23 ? plru1_39 : _GEN_2350; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2546 = _T_23 ? plru1_40 : _GEN_2351; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2547 = _T_23 ? plru1_41 : _GEN_2352; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2548 = _T_23 ? plru1_42 : _GEN_2353; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2549 = _T_23 ? plru1_43 : _GEN_2354; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2550 = _T_23 ? plru1_44 : _GEN_2355; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2551 = _T_23 ? plru1_45 : _GEN_2356; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2552 = _T_23 ? plru1_46 : _GEN_2357; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2553 = _T_23 ? plru1_47 : _GEN_2358; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2554 = _T_23 ? plru1_48 : _GEN_2359; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2555 = _T_23 ? plru1_49 : _GEN_2360; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2556 = _T_23 ? plru1_50 : _GEN_2361; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2557 = _T_23 ? plru1_51 : _GEN_2362; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2558 = _T_23 ? plru1_52 : _GEN_2363; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2559 = _T_23 ? plru1_53 : _GEN_2364; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2560 = _T_23 ? plru1_54 : _GEN_2365; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2561 = _T_23 ? plru1_55 : _GEN_2366; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2562 = _T_23 ? plru1_56 : _GEN_2367; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2563 = _T_23 ? plru1_57 : _GEN_2368; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2564 = _T_23 ? plru1_58 : _GEN_2369; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2565 = _T_23 ? plru1_59 : _GEN_2370; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2566 = _T_23 ? plru1_60 : _GEN_2371; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2567 = _T_23 ? plru1_61 : _GEN_2372; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2568 = _T_23 ? plru1_62 : _GEN_2373; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2569 = _T_23 ? plru1_63 : _GEN_2374; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2570 = _T_23 ? plru2_0 : _GEN_2375; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2571 = _T_23 ? plru2_1 : _GEN_2376; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2572 = _T_23 ? plru2_2 : _GEN_2377; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2573 = _T_23 ? plru2_3 : _GEN_2378; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2574 = _T_23 ? plru2_4 : _GEN_2379; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2575 = _T_23 ? plru2_5 : _GEN_2380; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2576 = _T_23 ? plru2_6 : _GEN_2381; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2577 = _T_23 ? plru2_7 : _GEN_2382; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2578 = _T_23 ? plru2_8 : _GEN_2383; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2579 = _T_23 ? plru2_9 : _GEN_2384; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2580 = _T_23 ? plru2_10 : _GEN_2385; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2581 = _T_23 ? plru2_11 : _GEN_2386; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2582 = _T_23 ? plru2_12 : _GEN_2387; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2583 = _T_23 ? plru2_13 : _GEN_2388; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2584 = _T_23 ? plru2_14 : _GEN_2389; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2585 = _T_23 ? plru2_15 : _GEN_2390; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2586 = _T_23 ? plru2_16 : _GEN_2391; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2587 = _T_23 ? plru2_17 : _GEN_2392; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2588 = _T_23 ? plru2_18 : _GEN_2393; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2589 = _T_23 ? plru2_19 : _GEN_2394; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2590 = _T_23 ? plru2_20 : _GEN_2395; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2591 = _T_23 ? plru2_21 : _GEN_2396; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2592 = _T_23 ? plru2_22 : _GEN_2397; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2593 = _T_23 ? plru2_23 : _GEN_2398; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2594 = _T_23 ? plru2_24 : _GEN_2399; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2595 = _T_23 ? plru2_25 : _GEN_2400; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2596 = _T_23 ? plru2_26 : _GEN_2401; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2597 = _T_23 ? plru2_27 : _GEN_2402; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2598 = _T_23 ? plru2_28 : _GEN_2403; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2599 = _T_23 ? plru2_29 : _GEN_2404; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2600 = _T_23 ? plru2_30 : _GEN_2405; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2601 = _T_23 ? plru2_31 : _GEN_2406; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2602 = _T_23 ? plru2_32 : _GEN_2407; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2603 = _T_23 ? plru2_33 : _GEN_2408; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2604 = _T_23 ? plru2_34 : _GEN_2409; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2605 = _T_23 ? plru2_35 : _GEN_2410; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2606 = _T_23 ? plru2_36 : _GEN_2411; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2607 = _T_23 ? plru2_37 : _GEN_2412; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2608 = _T_23 ? plru2_38 : _GEN_2413; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2609 = _T_23 ? plru2_39 : _GEN_2414; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2610 = _T_23 ? plru2_40 : _GEN_2415; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2611 = _T_23 ? plru2_41 : _GEN_2416; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2612 = _T_23 ? plru2_42 : _GEN_2417; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2613 = _T_23 ? plru2_43 : _GEN_2418; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2614 = _T_23 ? plru2_44 : _GEN_2419; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2615 = _T_23 ? plru2_45 : _GEN_2420; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2616 = _T_23 ? plru2_46 : _GEN_2421; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2617 = _T_23 ? plru2_47 : _GEN_2422; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2618 = _T_23 ? plru2_48 : _GEN_2423; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2619 = _T_23 ? plru2_49 : _GEN_2424; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2620 = _T_23 ? plru2_50 : _GEN_2425; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2621 = _T_23 ? plru2_51 : _GEN_2426; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2622 = _T_23 ? plru2_52 : _GEN_2427; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2623 = _T_23 ? plru2_53 : _GEN_2428; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2624 = _T_23 ? plru2_54 : _GEN_2429; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2625 = _T_23 ? plru2_55 : _GEN_2430; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2626 = _T_23 ? plru2_56 : _GEN_2431; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2627 = _T_23 ? plru2_57 : _GEN_2432; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2628 = _T_23 ? plru2_58 : _GEN_2433; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2629 = _T_23 ? plru2_59 : _GEN_2434; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2630 = _T_23 ? plru2_60 : _GEN_2435; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2631 = _T_23 ? plru2_61 : _GEN_2436; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2632 = _T_23 ? plru2_62 : _GEN_2437; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2633 = _T_23 ? plru2_63 : _GEN_2438; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire [63:0] _GEN_2634 = _T_23 ? 64'h0 : _GEN_2439; // @[Conditional.scala 39:67 Cache.scala 277:22]
  wire  _GEN_2635 = _T_16 ? _GEN_992 : fi_ready; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2637 = _T_16 ? _GEN_994 : _GEN_3; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2638 = _T_16 ? _GEN_995 : 128'h0; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_2639 = _T_16 ? _GEN_996 : 21'h0; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_2641 = _T_16 ? _GEN_999 : fi_ready; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2643 = _T_16 ? _GEN_1001 : _GEN_3; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2644 = _T_16 ? _GEN_1002 : 128'h0; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_2645 = _T_16 ? _GEN_1003 : 21'h0; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_2647 = _T_16 ? _GEN_1006 : fi_ready; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2649 = _T_16 ? _GEN_1008 : _GEN_3; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2650 = _T_16 ? _GEN_1009 : 128'h0; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_2651 = _T_16 ? _GEN_1010 : 21'h0; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_2653 = _T_16 ? _GEN_1013 : fi_ready; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2655 = _T_16 ? _GEN_1015 : _GEN_3; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2656 = _T_16 ? _GEN_1016 : 128'h0; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_2657 = _T_16 ? _GEN_1017 : 21'h0; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire [3:0] _GEN_2659 = _T_16 ? _GEN_1339 : _GEN_2440; // @[Conditional.scala 39:67]
  wire  _GEN_2660 = _T_16 ? _GEN_1340 : _GEN_2442; // @[Conditional.scala 39:67]
  wire  _GEN_2661 = _T_16 ? _GEN_1341 : _GEN_2443; // @[Conditional.scala 39:67]
  wire  _GEN_2662 = _T_16 ? _GEN_1342 : _GEN_2444; // @[Conditional.scala 39:67]
  wire  _GEN_2663 = _T_16 ? _GEN_1343 : _GEN_2445; // @[Conditional.scala 39:67]
  wire  _GEN_2664 = _T_16 ? _GEN_1344 : _GEN_2446; // @[Conditional.scala 39:67]
  wire  _GEN_2665 = _T_16 ? _GEN_1345 : _GEN_2447; // @[Conditional.scala 39:67]
  wire  _GEN_2666 = _T_16 ? _GEN_1346 : _GEN_2448; // @[Conditional.scala 39:67]
  wire  _GEN_2667 = _T_16 ? _GEN_1347 : _GEN_2449; // @[Conditional.scala 39:67]
  wire  _GEN_2668 = _T_16 ? _GEN_1348 : _GEN_2450; // @[Conditional.scala 39:67]
  wire  _GEN_2669 = _T_16 ? _GEN_1349 : _GEN_2451; // @[Conditional.scala 39:67]
  wire  _GEN_2670 = _T_16 ? _GEN_1350 : _GEN_2452; // @[Conditional.scala 39:67]
  wire  _GEN_2671 = _T_16 ? _GEN_1351 : _GEN_2453; // @[Conditional.scala 39:67]
  wire  _GEN_2672 = _T_16 ? _GEN_1352 : _GEN_2454; // @[Conditional.scala 39:67]
  wire  _GEN_2673 = _T_16 ? _GEN_1353 : _GEN_2455; // @[Conditional.scala 39:67]
  wire  _GEN_2674 = _T_16 ? _GEN_1354 : _GEN_2456; // @[Conditional.scala 39:67]
  wire  _GEN_2675 = _T_16 ? _GEN_1355 : _GEN_2457; // @[Conditional.scala 39:67]
  wire  _GEN_2676 = _T_16 ? _GEN_1356 : _GEN_2458; // @[Conditional.scala 39:67]
  wire  _GEN_2677 = _T_16 ? _GEN_1357 : _GEN_2459; // @[Conditional.scala 39:67]
  wire  _GEN_2678 = _T_16 ? _GEN_1358 : _GEN_2460; // @[Conditional.scala 39:67]
  wire  _GEN_2679 = _T_16 ? _GEN_1359 : _GEN_2461; // @[Conditional.scala 39:67]
  wire  _GEN_2680 = _T_16 ? _GEN_1360 : _GEN_2462; // @[Conditional.scala 39:67]
  wire  _GEN_2681 = _T_16 ? _GEN_1361 : _GEN_2463; // @[Conditional.scala 39:67]
  wire  _GEN_2682 = _T_16 ? _GEN_1362 : _GEN_2464; // @[Conditional.scala 39:67]
  wire  _GEN_2683 = _T_16 ? _GEN_1363 : _GEN_2465; // @[Conditional.scala 39:67]
  wire  _GEN_2684 = _T_16 ? _GEN_1364 : _GEN_2466; // @[Conditional.scala 39:67]
  wire  _GEN_2685 = _T_16 ? _GEN_1365 : _GEN_2467; // @[Conditional.scala 39:67]
  wire  _GEN_2686 = _T_16 ? _GEN_1366 : _GEN_2468; // @[Conditional.scala 39:67]
  wire  _GEN_2687 = _T_16 ? _GEN_1367 : _GEN_2469; // @[Conditional.scala 39:67]
  wire  _GEN_2688 = _T_16 ? _GEN_1368 : _GEN_2470; // @[Conditional.scala 39:67]
  wire  _GEN_2689 = _T_16 ? _GEN_1369 : _GEN_2471; // @[Conditional.scala 39:67]
  wire  _GEN_2690 = _T_16 ? _GEN_1370 : _GEN_2472; // @[Conditional.scala 39:67]
  wire  _GEN_2691 = _T_16 ? _GEN_1371 : _GEN_2473; // @[Conditional.scala 39:67]
  wire  _GEN_2692 = _T_16 ? _GEN_1372 : _GEN_2474; // @[Conditional.scala 39:67]
  wire  _GEN_2693 = _T_16 ? _GEN_1373 : _GEN_2475; // @[Conditional.scala 39:67]
  wire  _GEN_2694 = _T_16 ? _GEN_1374 : _GEN_2476; // @[Conditional.scala 39:67]
  wire  _GEN_2695 = _T_16 ? _GEN_1375 : _GEN_2477; // @[Conditional.scala 39:67]
  wire  _GEN_2696 = _T_16 ? _GEN_1376 : _GEN_2478; // @[Conditional.scala 39:67]
  wire  _GEN_2697 = _T_16 ? _GEN_1377 : _GEN_2479; // @[Conditional.scala 39:67]
  wire  _GEN_2698 = _T_16 ? _GEN_1378 : _GEN_2480; // @[Conditional.scala 39:67]
  wire  _GEN_2699 = _T_16 ? _GEN_1379 : _GEN_2481; // @[Conditional.scala 39:67]
  wire  _GEN_2700 = _T_16 ? _GEN_1380 : _GEN_2482; // @[Conditional.scala 39:67]
  wire  _GEN_2701 = _T_16 ? _GEN_1381 : _GEN_2483; // @[Conditional.scala 39:67]
  wire  _GEN_2702 = _T_16 ? _GEN_1382 : _GEN_2484; // @[Conditional.scala 39:67]
  wire  _GEN_2703 = _T_16 ? _GEN_1383 : _GEN_2485; // @[Conditional.scala 39:67]
  wire  _GEN_2704 = _T_16 ? _GEN_1384 : _GEN_2486; // @[Conditional.scala 39:67]
  wire  _GEN_2705 = _T_16 ? _GEN_1385 : _GEN_2487; // @[Conditional.scala 39:67]
  wire  _GEN_2706 = _T_16 ? _GEN_1386 : _GEN_2488; // @[Conditional.scala 39:67]
  wire  _GEN_2707 = _T_16 ? _GEN_1387 : _GEN_2489; // @[Conditional.scala 39:67]
  wire  _GEN_2708 = _T_16 ? _GEN_1388 : _GEN_2490; // @[Conditional.scala 39:67]
  wire  _GEN_2709 = _T_16 ? _GEN_1389 : _GEN_2491; // @[Conditional.scala 39:67]
  wire  _GEN_2710 = _T_16 ? _GEN_1390 : _GEN_2492; // @[Conditional.scala 39:67]
  wire  _GEN_2711 = _T_16 ? _GEN_1391 : _GEN_2493; // @[Conditional.scala 39:67]
  wire  _GEN_2712 = _T_16 ? _GEN_1392 : _GEN_2494; // @[Conditional.scala 39:67]
  wire  _GEN_2713 = _T_16 ? _GEN_1393 : _GEN_2495; // @[Conditional.scala 39:67]
  wire  _GEN_2714 = _T_16 ? _GEN_1394 : _GEN_2496; // @[Conditional.scala 39:67]
  wire  _GEN_2715 = _T_16 ? _GEN_1395 : _GEN_2497; // @[Conditional.scala 39:67]
  wire  _GEN_2716 = _T_16 ? _GEN_1396 : _GEN_2498; // @[Conditional.scala 39:67]
  wire  _GEN_2717 = _T_16 ? _GEN_1397 : _GEN_2499; // @[Conditional.scala 39:67]
  wire  _GEN_2718 = _T_16 ? _GEN_1398 : _GEN_2500; // @[Conditional.scala 39:67]
  wire  _GEN_2719 = _T_16 ? _GEN_1399 : _GEN_2501; // @[Conditional.scala 39:67]
  wire  _GEN_2720 = _T_16 ? _GEN_1400 : _GEN_2502; // @[Conditional.scala 39:67]
  wire  _GEN_2721 = _T_16 ? _GEN_1401 : _GEN_2503; // @[Conditional.scala 39:67]
  wire  _GEN_2722 = _T_16 ? _GEN_1402 : _GEN_2504; // @[Conditional.scala 39:67]
  wire  _GEN_2723 = _T_16 ? _GEN_1403 : _GEN_2505; // @[Conditional.scala 39:67]
  wire  _GEN_2724 = _T_16 ? _GEN_1404 : _GEN_2506; // @[Conditional.scala 39:67]
  wire  _GEN_2725 = _T_16 ? _GEN_1405 : _GEN_2507; // @[Conditional.scala 39:67]
  wire  _GEN_2726 = _T_16 ? _GEN_1406 : _GEN_2508; // @[Conditional.scala 39:67]
  wire  _GEN_2727 = _T_16 ? _GEN_1407 : _GEN_2509; // @[Conditional.scala 39:67]
  wire  _GEN_2728 = _T_16 ? _GEN_1408 : _GEN_2510; // @[Conditional.scala 39:67]
  wire  _GEN_2729 = _T_16 ? _GEN_1409 : _GEN_2511; // @[Conditional.scala 39:67]
  wire  _GEN_2730 = _T_16 ? _GEN_1410 : _GEN_2512; // @[Conditional.scala 39:67]
  wire  _GEN_2731 = _T_16 ? _GEN_1411 : _GEN_2513; // @[Conditional.scala 39:67]
  wire  _GEN_2732 = _T_16 ? _GEN_1412 : _GEN_2514; // @[Conditional.scala 39:67]
  wire  _GEN_2733 = _T_16 ? _GEN_1413 : _GEN_2515; // @[Conditional.scala 39:67]
  wire  _GEN_2734 = _T_16 ? _GEN_1414 : _GEN_2516; // @[Conditional.scala 39:67]
  wire  _GEN_2735 = _T_16 ? _GEN_1415 : _GEN_2517; // @[Conditional.scala 39:67]
  wire  _GEN_2736 = _T_16 ? _GEN_1416 : _GEN_2518; // @[Conditional.scala 39:67]
  wire  _GEN_2737 = _T_16 ? _GEN_1417 : _GEN_2519; // @[Conditional.scala 39:67]
  wire  _GEN_2738 = _T_16 ? _GEN_1418 : _GEN_2520; // @[Conditional.scala 39:67]
  wire  _GEN_2739 = _T_16 ? _GEN_1419 : _GEN_2521; // @[Conditional.scala 39:67]
  wire  _GEN_2740 = _T_16 ? _GEN_1420 : _GEN_2522; // @[Conditional.scala 39:67]
  wire  _GEN_2741 = _T_16 ? _GEN_1421 : _GEN_2523; // @[Conditional.scala 39:67]
  wire  _GEN_2742 = _T_16 ? _GEN_1422 : _GEN_2524; // @[Conditional.scala 39:67]
  wire  _GEN_2743 = _T_16 ? _GEN_1423 : _GEN_2525; // @[Conditional.scala 39:67]
  wire  _GEN_2744 = _T_16 ? _GEN_1424 : _GEN_2526; // @[Conditional.scala 39:67]
  wire  _GEN_2745 = _T_16 ? _GEN_1425 : _GEN_2527; // @[Conditional.scala 39:67]
  wire  _GEN_2746 = _T_16 ? _GEN_1426 : _GEN_2528; // @[Conditional.scala 39:67]
  wire  _GEN_2747 = _T_16 ? _GEN_1427 : _GEN_2529; // @[Conditional.scala 39:67]
  wire  _GEN_2748 = _T_16 ? _GEN_1428 : _GEN_2530; // @[Conditional.scala 39:67]
  wire  _GEN_2749 = _T_16 ? _GEN_1429 : _GEN_2531; // @[Conditional.scala 39:67]
  wire  _GEN_2750 = _T_16 ? _GEN_1430 : _GEN_2532; // @[Conditional.scala 39:67]
  wire  _GEN_2751 = _T_16 ? _GEN_1431 : _GEN_2533; // @[Conditional.scala 39:67]
  wire  _GEN_2752 = _T_16 ? _GEN_1432 : _GEN_2534; // @[Conditional.scala 39:67]
  wire  _GEN_2753 = _T_16 ? _GEN_1433 : _GEN_2535; // @[Conditional.scala 39:67]
  wire  _GEN_2754 = _T_16 ? _GEN_1434 : _GEN_2536; // @[Conditional.scala 39:67]
  wire  _GEN_2755 = _T_16 ? _GEN_1435 : _GEN_2537; // @[Conditional.scala 39:67]
  wire  _GEN_2756 = _T_16 ? _GEN_1436 : _GEN_2538; // @[Conditional.scala 39:67]
  wire  _GEN_2757 = _T_16 ? _GEN_1437 : _GEN_2539; // @[Conditional.scala 39:67]
  wire  _GEN_2758 = _T_16 ? _GEN_1438 : _GEN_2540; // @[Conditional.scala 39:67]
  wire  _GEN_2759 = _T_16 ? _GEN_1439 : _GEN_2541; // @[Conditional.scala 39:67]
  wire  _GEN_2760 = _T_16 ? _GEN_1440 : _GEN_2542; // @[Conditional.scala 39:67]
  wire  _GEN_2761 = _T_16 ? _GEN_1441 : _GEN_2543; // @[Conditional.scala 39:67]
  wire  _GEN_2762 = _T_16 ? _GEN_1442 : _GEN_2544; // @[Conditional.scala 39:67]
  wire  _GEN_2763 = _T_16 ? _GEN_1443 : _GEN_2545; // @[Conditional.scala 39:67]
  wire  _GEN_2764 = _T_16 ? _GEN_1444 : _GEN_2546; // @[Conditional.scala 39:67]
  wire  _GEN_2765 = _T_16 ? _GEN_1445 : _GEN_2547; // @[Conditional.scala 39:67]
  wire  _GEN_2766 = _T_16 ? _GEN_1446 : _GEN_2548; // @[Conditional.scala 39:67]
  wire  _GEN_2767 = _T_16 ? _GEN_1447 : _GEN_2549; // @[Conditional.scala 39:67]
  wire  _GEN_2768 = _T_16 ? _GEN_1448 : _GEN_2550; // @[Conditional.scala 39:67]
  wire  _GEN_2769 = _T_16 ? _GEN_1449 : _GEN_2551; // @[Conditional.scala 39:67]
  wire  _GEN_2770 = _T_16 ? _GEN_1450 : _GEN_2552; // @[Conditional.scala 39:67]
  wire  _GEN_2771 = _T_16 ? _GEN_1451 : _GEN_2553; // @[Conditional.scala 39:67]
  wire  _GEN_2772 = _T_16 ? _GEN_1452 : _GEN_2554; // @[Conditional.scala 39:67]
  wire  _GEN_2773 = _T_16 ? _GEN_1453 : _GEN_2555; // @[Conditional.scala 39:67]
  wire  _GEN_2774 = _T_16 ? _GEN_1454 : _GEN_2556; // @[Conditional.scala 39:67]
  wire  _GEN_2775 = _T_16 ? _GEN_1455 : _GEN_2557; // @[Conditional.scala 39:67]
  wire  _GEN_2776 = _T_16 ? _GEN_1456 : _GEN_2558; // @[Conditional.scala 39:67]
  wire  _GEN_2777 = _T_16 ? _GEN_1457 : _GEN_2559; // @[Conditional.scala 39:67]
  wire  _GEN_2778 = _T_16 ? _GEN_1458 : _GEN_2560; // @[Conditional.scala 39:67]
  wire  _GEN_2779 = _T_16 ? _GEN_1459 : _GEN_2561; // @[Conditional.scala 39:67]
  wire  _GEN_2780 = _T_16 ? _GEN_1460 : _GEN_2562; // @[Conditional.scala 39:67]
  wire  _GEN_2781 = _T_16 ? _GEN_1461 : _GEN_2563; // @[Conditional.scala 39:67]
  wire  _GEN_2782 = _T_16 ? _GEN_1462 : _GEN_2564; // @[Conditional.scala 39:67]
  wire  _GEN_2783 = _T_16 ? _GEN_1463 : _GEN_2565; // @[Conditional.scala 39:67]
  wire  _GEN_2784 = _T_16 ? _GEN_1464 : _GEN_2566; // @[Conditional.scala 39:67]
  wire  _GEN_2785 = _T_16 ? _GEN_1465 : _GEN_2567; // @[Conditional.scala 39:67]
  wire  _GEN_2786 = _T_16 ? _GEN_1466 : _GEN_2568; // @[Conditional.scala 39:67]
  wire  _GEN_2787 = _T_16 ? _GEN_1467 : _GEN_2569; // @[Conditional.scala 39:67]
  wire  _GEN_2788 = _T_16 ? _GEN_1468 : _GEN_2570; // @[Conditional.scala 39:67]
  wire  _GEN_2789 = _T_16 ? _GEN_1469 : _GEN_2571; // @[Conditional.scala 39:67]
  wire  _GEN_2790 = _T_16 ? _GEN_1470 : _GEN_2572; // @[Conditional.scala 39:67]
  wire  _GEN_2791 = _T_16 ? _GEN_1471 : _GEN_2573; // @[Conditional.scala 39:67]
  wire  _GEN_2792 = _T_16 ? _GEN_1472 : _GEN_2574; // @[Conditional.scala 39:67]
  wire  _GEN_2793 = _T_16 ? _GEN_1473 : _GEN_2575; // @[Conditional.scala 39:67]
  wire  _GEN_2794 = _T_16 ? _GEN_1474 : _GEN_2576; // @[Conditional.scala 39:67]
  wire  _GEN_2795 = _T_16 ? _GEN_1475 : _GEN_2577; // @[Conditional.scala 39:67]
  wire  _GEN_2796 = _T_16 ? _GEN_1476 : _GEN_2578; // @[Conditional.scala 39:67]
  wire  _GEN_2797 = _T_16 ? _GEN_1477 : _GEN_2579; // @[Conditional.scala 39:67]
  wire  _GEN_2798 = _T_16 ? _GEN_1478 : _GEN_2580; // @[Conditional.scala 39:67]
  wire  _GEN_2799 = _T_16 ? _GEN_1479 : _GEN_2581; // @[Conditional.scala 39:67]
  wire  _GEN_2800 = _T_16 ? _GEN_1480 : _GEN_2582; // @[Conditional.scala 39:67]
  wire  _GEN_2801 = _T_16 ? _GEN_1481 : _GEN_2583; // @[Conditional.scala 39:67]
  wire  _GEN_2802 = _T_16 ? _GEN_1482 : _GEN_2584; // @[Conditional.scala 39:67]
  wire  _GEN_2803 = _T_16 ? _GEN_1483 : _GEN_2585; // @[Conditional.scala 39:67]
  wire  _GEN_2804 = _T_16 ? _GEN_1484 : _GEN_2586; // @[Conditional.scala 39:67]
  wire  _GEN_2805 = _T_16 ? _GEN_1485 : _GEN_2587; // @[Conditional.scala 39:67]
  wire  _GEN_2806 = _T_16 ? _GEN_1486 : _GEN_2588; // @[Conditional.scala 39:67]
  wire  _GEN_2807 = _T_16 ? _GEN_1487 : _GEN_2589; // @[Conditional.scala 39:67]
  wire  _GEN_2808 = _T_16 ? _GEN_1488 : _GEN_2590; // @[Conditional.scala 39:67]
  wire  _GEN_2809 = _T_16 ? _GEN_1489 : _GEN_2591; // @[Conditional.scala 39:67]
  wire  _GEN_2810 = _T_16 ? _GEN_1490 : _GEN_2592; // @[Conditional.scala 39:67]
  wire  _GEN_2811 = _T_16 ? _GEN_1491 : _GEN_2593; // @[Conditional.scala 39:67]
  wire  _GEN_2812 = _T_16 ? _GEN_1492 : _GEN_2594; // @[Conditional.scala 39:67]
  wire  _GEN_2813 = _T_16 ? _GEN_1493 : _GEN_2595; // @[Conditional.scala 39:67]
  wire  _GEN_2814 = _T_16 ? _GEN_1494 : _GEN_2596; // @[Conditional.scala 39:67]
  wire  _GEN_2815 = _T_16 ? _GEN_1495 : _GEN_2597; // @[Conditional.scala 39:67]
  wire  _GEN_2816 = _T_16 ? _GEN_1496 : _GEN_2598; // @[Conditional.scala 39:67]
  wire  _GEN_2817 = _T_16 ? _GEN_1497 : _GEN_2599; // @[Conditional.scala 39:67]
  wire  _GEN_2818 = _T_16 ? _GEN_1498 : _GEN_2600; // @[Conditional.scala 39:67]
  wire  _GEN_2819 = _T_16 ? _GEN_1499 : _GEN_2601; // @[Conditional.scala 39:67]
  wire  _GEN_2820 = _T_16 ? _GEN_1500 : _GEN_2602; // @[Conditional.scala 39:67]
  wire  _GEN_2821 = _T_16 ? _GEN_1501 : _GEN_2603; // @[Conditional.scala 39:67]
  wire  _GEN_2822 = _T_16 ? _GEN_1502 : _GEN_2604; // @[Conditional.scala 39:67]
  wire  _GEN_2823 = _T_16 ? _GEN_1503 : _GEN_2605; // @[Conditional.scala 39:67]
  wire  _GEN_2824 = _T_16 ? _GEN_1504 : _GEN_2606; // @[Conditional.scala 39:67]
  wire  _GEN_2825 = _T_16 ? _GEN_1505 : _GEN_2607; // @[Conditional.scala 39:67]
  wire  _GEN_2826 = _T_16 ? _GEN_1506 : _GEN_2608; // @[Conditional.scala 39:67]
  wire  _GEN_2827 = _T_16 ? _GEN_1507 : _GEN_2609; // @[Conditional.scala 39:67]
  wire  _GEN_2828 = _T_16 ? _GEN_1508 : _GEN_2610; // @[Conditional.scala 39:67]
  wire  _GEN_2829 = _T_16 ? _GEN_1509 : _GEN_2611; // @[Conditional.scala 39:67]
  wire  _GEN_2830 = _T_16 ? _GEN_1510 : _GEN_2612; // @[Conditional.scala 39:67]
  wire  _GEN_2831 = _T_16 ? _GEN_1511 : _GEN_2613; // @[Conditional.scala 39:67]
  wire  _GEN_2832 = _T_16 ? _GEN_1512 : _GEN_2614; // @[Conditional.scala 39:67]
  wire  _GEN_2833 = _T_16 ? _GEN_1513 : _GEN_2615; // @[Conditional.scala 39:67]
  wire  _GEN_2834 = _T_16 ? _GEN_1514 : _GEN_2616; // @[Conditional.scala 39:67]
  wire  _GEN_2835 = _T_16 ? _GEN_1515 : _GEN_2617; // @[Conditional.scala 39:67]
  wire  _GEN_2836 = _T_16 ? _GEN_1516 : _GEN_2618; // @[Conditional.scala 39:67]
  wire  _GEN_2837 = _T_16 ? _GEN_1517 : _GEN_2619; // @[Conditional.scala 39:67]
  wire  _GEN_2838 = _T_16 ? _GEN_1518 : _GEN_2620; // @[Conditional.scala 39:67]
  wire  _GEN_2839 = _T_16 ? _GEN_1519 : _GEN_2621; // @[Conditional.scala 39:67]
  wire  _GEN_2840 = _T_16 ? _GEN_1520 : _GEN_2622; // @[Conditional.scala 39:67]
  wire  _GEN_2841 = _T_16 ? _GEN_1521 : _GEN_2623; // @[Conditional.scala 39:67]
  wire  _GEN_2842 = _T_16 ? _GEN_1522 : _GEN_2624; // @[Conditional.scala 39:67]
  wire  _GEN_2843 = _T_16 ? _GEN_1523 : _GEN_2625; // @[Conditional.scala 39:67]
  wire  _GEN_2844 = _T_16 ? _GEN_1524 : _GEN_2626; // @[Conditional.scala 39:67]
  wire  _GEN_2845 = _T_16 ? _GEN_1525 : _GEN_2627; // @[Conditional.scala 39:67]
  wire  _GEN_2846 = _T_16 ? _GEN_1526 : _GEN_2628; // @[Conditional.scala 39:67]
  wire  _GEN_2847 = _T_16 ? _GEN_1527 : _GEN_2629; // @[Conditional.scala 39:67]
  wire  _GEN_2848 = _T_16 ? _GEN_1528 : _GEN_2630; // @[Conditional.scala 39:67]
  wire  _GEN_2849 = _T_16 ? _GEN_1529 : _GEN_2631; // @[Conditional.scala 39:67]
  wire  _GEN_2850 = _T_16 ? _GEN_1530 : _GEN_2632; // @[Conditional.scala 39:67]
  wire  _GEN_2851 = _T_16 ? _GEN_1531 : _GEN_2633; // @[Conditional.scala 39:67]
  wire  _GEN_2852 = _T_16 ? _GEN_27 : _GEN_2441; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_2853 = _T_16 ? 64'h0 : _GEN_2634; // @[Conditional.scala 39:67 Cache.scala 277:22]
  wire [3:0] _GEN_2856 = _T_13 ? _GEN_990 : _GEN_2659; // @[Conditional.scala 39:67]
  wire  _GEN_2857 = _T_13 ? fi_ready : _GEN_2635; // @[Conditional.scala 39:67]
  wire  _GEN_2858 = _T_13 ? 1'h0 : _T_16 & _T_17; // @[Conditional.scala 39:67 Cache.scala 110:14]
  wire [5:0] _GEN_2859 = _T_13 ? _GEN_3 : _GEN_2637; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2860 = _T_13 ? 128'h0 : _GEN_2638; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_2861 = _T_13 ? 21'h0 : _GEN_2639; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_2862 = _T_13 ? 1'h0 : _T_16 & _GEN_997; // @[Conditional.scala 39:67 Cache.scala 118:18]
  wire  _GEN_2863 = _T_13 ? fi_ready : _GEN_2641; // @[Conditional.scala 39:67]
  wire  _GEN_2864 = _T_13 ? 1'h0 : _T_16 & _T_18; // @[Conditional.scala 39:67 Cache.scala 110:14]
  wire [5:0] _GEN_2865 = _T_13 ? _GEN_3 : _GEN_2643; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2866 = _T_13 ? 128'h0 : _GEN_2644; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_2867 = _T_13 ? 21'h0 : _GEN_2645; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_2868 = _T_13 ? 1'h0 : _T_16 & _GEN_1004; // @[Conditional.scala 39:67 Cache.scala 118:18]
  wire  _GEN_2869 = _T_13 ? fi_ready : _GEN_2647; // @[Conditional.scala 39:67]
  wire  _GEN_2870 = _T_13 ? 1'h0 : _T_16 & _T_19; // @[Conditional.scala 39:67 Cache.scala 110:14]
  wire [5:0] _GEN_2871 = _T_13 ? _GEN_3 : _GEN_2649; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2872 = _T_13 ? 128'h0 : _GEN_2650; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_2873 = _T_13 ? 21'h0 : _GEN_2651; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_2874 = _T_13 ? 1'h0 : _T_16 & _GEN_1011; // @[Conditional.scala 39:67 Cache.scala 118:18]
  wire  _GEN_2875 = _T_13 ? fi_ready : _GEN_2653; // @[Conditional.scala 39:67]
  wire  _GEN_2876 = _T_13 ? 1'h0 : _T_16 & _T_20; // @[Conditional.scala 39:67 Cache.scala 110:14]
  wire [5:0] _GEN_2877 = _T_13 ? _GEN_3 : _GEN_2655; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2878 = _T_13 ? 128'h0 : _GEN_2656; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_2879 = _T_13 ? 21'h0 : _GEN_2657; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_2880 = _T_13 ? 1'h0 : _T_16 & _GEN_1018; // @[Conditional.scala 39:67 Cache.scala 118:18]
  wire [63:0] _GEN_3074 = _T_13 ? 64'h0 : _GEN_2853; // @[Conditional.scala 39:67 Cache.scala 277:22]
  wire [3:0] _GEN_3075 = _T_11 ? _GEN_984 : _GEN_2856; // @[Conditional.scala 39:67]
  wire  _GEN_3078 = _T_11 ? fi_ready : _GEN_2857; // @[Conditional.scala 39:67]
  wire  _GEN_3079 = _T_11 ? 1'h0 : _GEN_2858; // @[Conditional.scala 39:67 Cache.scala 110:14]
  wire [5:0] _GEN_3080 = _T_11 ? _GEN_3 : _GEN_2859; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_3081 = _T_11 ? 128'h0 : _GEN_2860; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_3082 = _T_11 ? 21'h0 : _GEN_2861; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_3083 = _T_11 ? 1'h0 : _GEN_2862; // @[Conditional.scala 39:67 Cache.scala 118:18]
  wire  _GEN_3084 = _T_11 ? fi_ready : _GEN_2863; // @[Conditional.scala 39:67]
  wire  _GEN_3085 = _T_11 ? 1'h0 : _GEN_2864; // @[Conditional.scala 39:67 Cache.scala 110:14]
  wire [5:0] _GEN_3086 = _T_11 ? _GEN_3 : _GEN_2865; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_3087 = _T_11 ? 128'h0 : _GEN_2866; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_3088 = _T_11 ? 21'h0 : _GEN_2867; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_3089 = _T_11 ? 1'h0 : _GEN_2868; // @[Conditional.scala 39:67 Cache.scala 118:18]
  wire  _GEN_3090 = _T_11 ? fi_ready : _GEN_2869; // @[Conditional.scala 39:67]
  wire  _GEN_3091 = _T_11 ? 1'h0 : _GEN_2870; // @[Conditional.scala 39:67 Cache.scala 110:14]
  wire [5:0] _GEN_3092 = _T_11 ? _GEN_3 : _GEN_2871; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_3093 = _T_11 ? 128'h0 : _GEN_2872; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_3094 = _T_11 ? 21'h0 : _GEN_2873; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_3095 = _T_11 ? 1'h0 : _GEN_2874; // @[Conditional.scala 39:67 Cache.scala 118:18]
  wire  _GEN_3096 = _T_11 ? fi_ready : _GEN_2875; // @[Conditional.scala 39:67]
  wire  _GEN_3097 = _T_11 ? 1'h0 : _GEN_2876; // @[Conditional.scala 39:67 Cache.scala 110:14]
  wire [5:0] _GEN_3098 = _T_11 ? _GEN_3 : _GEN_2877; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_3099 = _T_11 ? 128'h0 : _GEN_2878; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_3100 = _T_11 ? 21'h0 : _GEN_2879; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_3101 = _T_11 ? 1'h0 : _GEN_2880; // @[Conditional.scala 39:67 Cache.scala 118:18]
  wire [63:0] _GEN_3295 = _T_11 ? 64'h0 : _GEN_3074; // @[Conditional.scala 39:67 Cache.scala 277:22]
  wire  _io_out_req_valid_T = state == 4'h1; // @[Cache.scala 504:27]
  wire  _io_out_req_valid_T_1 = state == 4'h4; // @[Cache.scala 505:27]
  wire  _io_out_req_valid_T_2 = state == 4'h1 | _io_out_req_valid_T_1; // @[Cache.scala 504:45]
  wire  _io_out_req_valid_T_3 = state == 4'h5; // @[Cache.scala 506:27]
  wire [27:0] io_out_req_bits_addr_hi = s2_addr[31:4]; // @[Cache.scala 512:37]
  wire [31:0] _io_out_req_bits_addr_T = {io_out_req_bits_addr_hi,4'h0}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_3534 = _io_out_req_valid_T ? _io_out_req_bits_addr_T : 32'h0; // @[Cache.scala 511:33 Cache.scala 512:23 Cache.scala 510:21]
  wire [31:0] _io_out_req_bits_addr_T_1 = {1'h1,s2_reg_tag_r,s2_idx,4'h0}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_3537 = _io_out_req_valid_T_1 ? s2_reg_dat_w[63:0] : 64'h0; // @[Cache.scala 527:34 Cache.scala 528:24 Cache.scala 526:22]
  wire  _io_out_resp_ready_T_1 = state == 4'h6; // @[Cache.scala 549:28]

  assign io_sram0_addr = sram_0_io_addr; 
  assign io_sram0_cen = ~sram_0_io_en; 
  assign io_sram0_wen = ~sram_0_io_wen; 
  assign io_sram0_wdata = sram_0_io_wdata; 
  assign io_sram1_addr = sram_1_io_addr; 
  assign io_sram1_cen = ~sram_1_io_en; 
  assign io_sram1_wen = ~sram_1_io_wen; 
  assign io_sram1_wdata = sram_1_io_wdata; 
  assign io_sram2_addr = sram_2_io_addr; 
  assign io_sram2_cen = ~sram_2_io_en; 
  assign io_sram2_wen = ~sram_2_io_wen; 
  assign io_sram2_wdata = sram_2_io_wdata; 
  assign io_sram3_addr = sram_3_io_addr; 
  assign io_sram3_cen = ~sram_3_io_en; 
  assign io_sram3_wen = ~sram_3_io_wen; 
  assign io_sram3_wdata = sram_3_io_wdata; 

  assign sram_0_io_rdata = io_sram0_rdata;
  assign sram_3_io_rdata = io_sram3_rdata;
  assign sram_2_io_rdata = io_sram2_rdata;
  assign sram_1_io_rdata = io_sram1_rdata;
/*
  ysyx_210340_Sram sram_0 ( // @[Cache.scala 91:22]
    .clock(sram_0_clock),
    .io_en(sram_0_io_en),
    .io_wen(sram_0_io_wen),
    .io_addr(sram_0_io_addr),
    .io_wdata(sram_0_io_wdata),
    .io_rdata(sram_0_io_rdata)
  );
  ysyx_210340_Sram sram_1 ( // @[Cache.scala 91:22]
    .clock(sram_1_clock),
    .io_en(sram_1_io_en),
    .io_wen(sram_1_io_wen),
    .io_addr(sram_1_io_addr),
    .io_wdata(sram_1_io_wdata),
    .io_rdata(sram_1_io_rdata)
  );
  ysyx_210340_Sram sram_2 ( // @[Cache.scala 91:22]
    .clock(sram_2_clock),
    .io_en(sram_2_io_en),
    .io_wen(sram_2_io_wen),
    .io_addr(sram_2_io_addr),
    .io_wdata(sram_2_io_wdata),
    .io_rdata(sram_2_io_rdata)
  );
  ysyx_210340_Sram sram_3 ( // @[Cache.scala 91:22]
    .clock(sram_3_clock),
    .io_en(sram_3_io_en),
    .io_wen(sram_3_io_wen),
    .io_addr(sram_3_io_addr),
    .io_wdata(sram_3_io_wdata),
    .io_rdata(sram_3_io_rdata)
  );
*/
  ysyx_210340_Meta meta_0 ( // @[Cache.scala 99:22]
    .clock(meta_0_clock),
    .reset(meta_0_reset),
    .io_idx(meta_0_io_idx),
    .io_tag_r(meta_0_io_tag_r),
    .io_tag_w(meta_0_io_tag_w),
    .io_tag_wen(meta_0_io_tag_wen),
    .io_dirty_r(meta_0_io_dirty_r),
    .io_dirty_w(meta_0_io_dirty_w),
    .io_dirty_wen(meta_0_io_dirty_wen),
    .io_valid_r(meta_0_io_valid_r),
    .io_invalidate(meta_0_io_invalidate),
    .io_dirty_r_async(meta_0_io_dirty_r_async),
    .io_valid_r_async(meta_0_io_valid_r_async)
  );
  ysyx_210340_Meta meta_1 ( // @[Cache.scala 99:22]
    .clock(meta_1_clock),
    .reset(meta_1_reset),
    .io_idx(meta_1_io_idx),
    .io_tag_r(meta_1_io_tag_r),
    .io_tag_w(meta_1_io_tag_w),
    .io_tag_wen(meta_1_io_tag_wen),
    .io_dirty_r(meta_1_io_dirty_r),
    .io_dirty_w(meta_1_io_dirty_w),
    .io_dirty_wen(meta_1_io_dirty_wen),
    .io_valid_r(meta_1_io_valid_r),
    .io_invalidate(meta_1_io_invalidate),
    .io_dirty_r_async(meta_1_io_dirty_r_async),
    .io_valid_r_async(meta_1_io_valid_r_async)
  );
  ysyx_210340_Meta meta_2 ( // @[Cache.scala 99:22]
    .clock(meta_2_clock),
    .reset(meta_2_reset),
    .io_idx(meta_2_io_idx),
    .io_tag_r(meta_2_io_tag_r),
    .io_tag_w(meta_2_io_tag_w),
    .io_tag_wen(meta_2_io_tag_wen),
    .io_dirty_r(meta_2_io_dirty_r),
    .io_dirty_w(meta_2_io_dirty_w),
    .io_dirty_wen(meta_2_io_dirty_wen),
    .io_valid_r(meta_2_io_valid_r),
    .io_invalidate(meta_2_io_invalidate),
    .io_dirty_r_async(meta_2_io_dirty_r_async),
    .io_valid_r_async(meta_2_io_valid_r_async)
  );
  ysyx_210340_Meta meta_3 ( // @[Cache.scala 99:22]
    .clock(meta_3_clock),
    .reset(meta_3_reset),
    .io_idx(meta_3_io_idx),
    .io_tag_r(meta_3_io_tag_r),
    .io_tag_w(meta_3_io_tag_w),
    .io_tag_wen(meta_3_io_tag_wen),
    .io_dirty_r(meta_3_io_dirty_r),
    .io_dirty_w(meta_3_io_dirty_w),
    .io_dirty_wen(meta_3_io_dirty_wen),
    .io_valid_r(meta_3_io_valid_r),
    .io_invalidate(meta_3_io_invalidate),
    .io_dirty_r_async(meta_3_io_dirty_r_async),
    .io_valid_r_async(meta_3_io_valid_r_async)
  );
  assign io_in_req_ready = fi_ready & ~fi_valid; // @[Cache.scala 275:34]
  assign io_in_resp_valid = s2_hit_real & ~s2_wen & state != 4'h8 | _hit_ready_T; // @[Cache.scala 276:71]
  assign io_in_resp_bits_rdata = _T_2 ? _GEN_228 : _GEN_3295; // @[Conditional.scala 40:58]
  assign io_out_req_valid = _io_out_req_valid_T_2 | _io_out_req_valid_T_3; // @[Cache.scala 505:46]
  assign io_out_req_bits_addr = _io_out_req_valid_T_1 ? _io_out_req_bits_addr_T_1 : _GEN_3534; // @[Cache.scala 514:34 Cache.scala 517:23]
  assign io_out_req_bits_aen = _io_out_req_valid_T | _io_out_req_valid_T_1; // @[Cache.scala 522:48]
  assign io_out_req_bits_ren = state == 4'h1; // @[Cache.scala 525:30]
  assign io_out_req_bits_wdata = _io_out_req_valid_T_3 ? s2_reg_dat_w[127:64] : _GEN_3537; // @[Cache.scala 530:34 Cache.scala 531:24]
  assign io_out_req_bits_wlast = state == 4'h5; // @[Cache.scala 540:32]
  assign io_out_req_bits_wen = _io_out_req_valid_T_1 | _io_out_req_valid_T_3; // @[Cache.scala 542:49]
  assign io_out_resp_ready = state == 4'h2 | _io_out_resp_ready_T_1; // @[Cache.scala 548:47]
  // assign sram_0_clock = clock;
  assign sram_0_io_en = _T_2 ? _GEN_967 : _GEN_3078; // @[Conditional.scala 40:58]
  assign sram_0_io_wen = _T_2 ? _GEN_968 : _GEN_3079; // @[Conditional.scala 40:58]
  assign sram_0_io_addr = _T_2 ? _GEN_969 : _GEN_3080; // @[Conditional.scala 40:58]
  assign sram_0_io_wdata = _T_2 ? _GEN_970 : _GEN_3081; // @[Conditional.scala 40:58]
  // assign sram_1_clock = clock;
  assign sram_1_io_en = _T_2 ? _GEN_971 : _GEN_3084; // @[Conditional.scala 40:58]
  assign sram_1_io_wen = _T_2 ? _GEN_972 : _GEN_3085; // @[Conditional.scala 40:58]
  assign sram_1_io_addr = _T_2 ? _GEN_973 : _GEN_3086; // @[Conditional.scala 40:58]
  assign sram_1_io_wdata = _T_2 ? _GEN_974 : _GEN_3087; // @[Conditional.scala 40:58]
  // assign sram_2_clock = clock;
  assign sram_2_io_en = _T_2 ? _GEN_975 : _GEN_3090; // @[Conditional.scala 40:58]
  assign sram_2_io_wen = _T_2 ? _GEN_976 : _GEN_3091; // @[Conditional.scala 40:58]
  assign sram_2_io_addr = _T_2 ? _GEN_977 : _GEN_3092; // @[Conditional.scala 40:58]
  assign sram_2_io_wdata = _T_2 ? _GEN_978 : _GEN_3093; // @[Conditional.scala 40:58]
  // assign sram_3_clock = clock;
  assign sram_3_io_en = _T_2 ? _GEN_979 : _GEN_3096; // @[Conditional.scala 40:58]
  assign sram_3_io_wen = _T_2 ? _GEN_980 : _GEN_3097; // @[Conditional.scala 40:58]
  assign sram_3_io_addr = _T_2 ? _GEN_981 : _GEN_3098; // @[Conditional.scala 40:58]
  assign sram_3_io_wdata = _T_2 ? _GEN_982 : _GEN_3099; // @[Conditional.scala 40:58]
  assign meta_0_clock = clock;
  assign meta_0_reset = reset;
  assign meta_0_io_idx = _T_2 ? _GEN_969 : _GEN_3080; // @[Conditional.scala 40:58]
  assign meta_0_io_tag_w = _T_2 ? 21'h0 : _GEN_3082; // @[Conditional.scala 40:58 Cache.scala 116:16]
  assign meta_0_io_tag_wen = _T_2 ? 1'h0 : _GEN_3079; // @[Conditional.scala 40:58 Cache.scala 117:18]
  assign meta_0_io_dirty_w = _T_2 ? _GEN_968 : _GEN_3083; // @[Conditional.scala 40:58]
  assign meta_0_io_dirty_wen = _T_2 ? _GEN_968 : _GEN_3079; // @[Conditional.scala 40:58]
  assign meta_0_io_invalidate = fi_valid & fi_ready; // @[Cache.scala 163:26]
  assign meta_1_clock = clock;
  assign meta_1_reset = reset;
  assign meta_1_io_idx = _T_2 ? _GEN_973 : _GEN_3086; // @[Conditional.scala 40:58]
  assign meta_1_io_tag_w = _T_2 ? 21'h0 : _GEN_3088; // @[Conditional.scala 40:58 Cache.scala 116:16]
  assign meta_1_io_tag_wen = _T_2 ? 1'h0 : _GEN_3085; // @[Conditional.scala 40:58 Cache.scala 117:18]
  assign meta_1_io_dirty_w = _T_2 ? _GEN_972 : _GEN_3089; // @[Conditional.scala 40:58]
  assign meta_1_io_dirty_wen = _T_2 ? _GEN_972 : _GEN_3085; // @[Conditional.scala 40:58]
  assign meta_1_io_invalidate = fi_valid & fi_ready; // @[Cache.scala 163:26]
  assign meta_2_clock = clock;
  assign meta_2_reset = reset;
  assign meta_2_io_idx = _T_2 ? _GEN_977 : _GEN_3092; // @[Conditional.scala 40:58]
  assign meta_2_io_tag_w = _T_2 ? 21'h0 : _GEN_3094; // @[Conditional.scala 40:58 Cache.scala 116:16]
  assign meta_2_io_tag_wen = _T_2 ? 1'h0 : _GEN_3091; // @[Conditional.scala 40:58 Cache.scala 117:18]
  assign meta_2_io_dirty_w = _T_2 ? _GEN_976 : _GEN_3095; // @[Conditional.scala 40:58]
  assign meta_2_io_dirty_wen = _T_2 ? _GEN_976 : _GEN_3091; // @[Conditional.scala 40:58]
  assign meta_2_io_invalidate = fi_valid & fi_ready; // @[Cache.scala 163:26]
  assign meta_3_clock = clock;
  assign meta_3_reset = reset;
  assign meta_3_io_idx = _T_2 ? _GEN_981 : _GEN_3098; // @[Conditional.scala 40:58]
  assign meta_3_io_tag_w = _T_2 ? 21'h0 : _GEN_3100; // @[Conditional.scala 40:58 Cache.scala 116:16]
  assign meta_3_io_tag_wen = _T_2 ? 1'h0 : _GEN_3097; // @[Conditional.scala 40:58 Cache.scala 117:18]
  assign meta_3_io_dirty_w = _T_2 ? _GEN_980 : _GEN_3101; // @[Conditional.scala 40:58]
  assign meta_3_io_dirty_wen = _T_2 ? _GEN_980 : _GEN_3097; // @[Conditional.scala 40:58]
  assign meta_3_io_invalidate = fi_valid & fi_ready; // @[Cache.scala 163:26]
  always @(posedge clock) begin
    if (reset) begin // @[Cache.scala 131:22]
      plru0_0 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_0 <= _GEN_229;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_0 <= _GEN_2660;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_1 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_1 <= _GEN_230;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_1 <= _GEN_2661;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_2 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_2 <= _GEN_231;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_2 <= _GEN_2662;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_3 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_3 <= _GEN_232;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_3 <= _GEN_2663;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_4 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_4 <= _GEN_233;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_4 <= _GEN_2664;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_5 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_5 <= _GEN_234;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_5 <= _GEN_2665;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_6 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_6 <= _GEN_235;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_6 <= _GEN_2666;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_7 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_7 <= _GEN_236;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_7 <= _GEN_2667;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_8 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_8 <= _GEN_237;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_8 <= _GEN_2668;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_9 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_9 <= _GEN_238;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_9 <= _GEN_2669;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_10 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_10 <= _GEN_239;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_10 <= _GEN_2670;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_11 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_11 <= _GEN_240;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_11 <= _GEN_2671;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_12 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_12 <= _GEN_241;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_12 <= _GEN_2672;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_13 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_13 <= _GEN_242;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_13 <= _GEN_2673;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_14 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_14 <= _GEN_243;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_14 <= _GEN_2674;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_15 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_15 <= _GEN_244;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_15 <= _GEN_2675;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_16 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_16 <= _GEN_245;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_16 <= _GEN_2676;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_17 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_17 <= _GEN_246;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_17 <= _GEN_2677;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_18 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_18 <= _GEN_247;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_18 <= _GEN_2678;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_19 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_19 <= _GEN_248;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_19 <= _GEN_2679;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_20 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_20 <= _GEN_249;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_20 <= _GEN_2680;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_21 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_21 <= _GEN_250;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_21 <= _GEN_2681;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_22 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_22 <= _GEN_251;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_22 <= _GEN_2682;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_23 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_23 <= _GEN_252;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_23 <= _GEN_2683;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_24 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_24 <= _GEN_253;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_24 <= _GEN_2684;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_25 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_25 <= _GEN_254;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_25 <= _GEN_2685;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_26 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_26 <= _GEN_255;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_26 <= _GEN_2686;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_27 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_27 <= _GEN_256;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_27 <= _GEN_2687;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_28 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_28 <= _GEN_257;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_28 <= _GEN_2688;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_29 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_29 <= _GEN_258;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_29 <= _GEN_2689;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_30 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_30 <= _GEN_259;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_30 <= _GEN_2690;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_31 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_31 <= _GEN_260;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_31 <= _GEN_2691;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_32 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_32 <= _GEN_261;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_32 <= _GEN_2692;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_33 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_33 <= _GEN_262;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_33 <= _GEN_2693;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_34 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_34 <= _GEN_263;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_34 <= _GEN_2694;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_35 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_35 <= _GEN_264;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_35 <= _GEN_2695;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_36 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_36 <= _GEN_265;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_36 <= _GEN_2696;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_37 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_37 <= _GEN_266;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_37 <= _GEN_2697;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_38 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_38 <= _GEN_267;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_38 <= _GEN_2698;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_39 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_39 <= _GEN_268;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_39 <= _GEN_2699;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_40 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_40 <= _GEN_269;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_40 <= _GEN_2700;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_41 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_41 <= _GEN_270;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_41 <= _GEN_2701;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_42 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_42 <= _GEN_271;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_42 <= _GEN_2702;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_43 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_43 <= _GEN_272;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_43 <= _GEN_2703;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_44 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_44 <= _GEN_273;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_44 <= _GEN_2704;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_45 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_45 <= _GEN_274;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_45 <= _GEN_2705;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_46 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_46 <= _GEN_275;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_46 <= _GEN_2706;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_47 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_47 <= _GEN_276;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_47 <= _GEN_2707;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_48 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_48 <= _GEN_277;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_48 <= _GEN_2708;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_49 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_49 <= _GEN_278;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_49 <= _GEN_2709;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_50 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_50 <= _GEN_279;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_50 <= _GEN_2710;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_51 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_51 <= _GEN_280;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_51 <= _GEN_2711;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_52 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_52 <= _GEN_281;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_52 <= _GEN_2712;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_53 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_53 <= _GEN_282;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_53 <= _GEN_2713;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_54 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_54 <= _GEN_283;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_54 <= _GEN_2714;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_55 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_55 <= _GEN_284;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_55 <= _GEN_2715;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_56 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_56 <= _GEN_285;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_56 <= _GEN_2716;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_57 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_57 <= _GEN_286;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_57 <= _GEN_2717;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_58 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_58 <= _GEN_287;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_58 <= _GEN_2718;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_59 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_59 <= _GEN_288;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_59 <= _GEN_2719;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_60 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_60 <= _GEN_289;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_60 <= _GEN_2720;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_61 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_61 <= _GEN_290;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_61 <= _GEN_2721;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_62 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_62 <= _GEN_291;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_62 <= _GEN_2722;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_63 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_63 <= _GEN_292;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_63 <= _GEN_2723;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_0 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_0 <= _GEN_421;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_0 <= _GEN_2724;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_1 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_1 <= _GEN_422;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_1 <= _GEN_2725;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_2 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_2 <= _GEN_423;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_2 <= _GEN_2726;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_3 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_3 <= _GEN_424;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_3 <= _GEN_2727;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_4 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_4 <= _GEN_425;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_4 <= _GEN_2728;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_5 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_5 <= _GEN_426;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_5 <= _GEN_2729;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_6 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_6 <= _GEN_427;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_6 <= _GEN_2730;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_7 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_7 <= _GEN_428;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_7 <= _GEN_2731;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_8 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_8 <= _GEN_429;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_8 <= _GEN_2732;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_9 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_9 <= _GEN_430;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_9 <= _GEN_2733;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_10 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_10 <= _GEN_431;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_10 <= _GEN_2734;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_11 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_11 <= _GEN_432;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_11 <= _GEN_2735;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_12 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_12 <= _GEN_433;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_12 <= _GEN_2736;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_13 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_13 <= _GEN_434;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_13 <= _GEN_2737;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_14 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_14 <= _GEN_435;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_14 <= _GEN_2738;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_15 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_15 <= _GEN_436;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_15 <= _GEN_2739;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_16 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_16 <= _GEN_437;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_16 <= _GEN_2740;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_17 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_17 <= _GEN_438;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_17 <= _GEN_2741;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_18 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_18 <= _GEN_439;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_18 <= _GEN_2742;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_19 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_19 <= _GEN_440;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_19 <= _GEN_2743;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_20 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_20 <= _GEN_441;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_20 <= _GEN_2744;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_21 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_21 <= _GEN_442;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_21 <= _GEN_2745;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_22 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_22 <= _GEN_443;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_22 <= _GEN_2746;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_23 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_23 <= _GEN_444;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_23 <= _GEN_2747;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_24 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_24 <= _GEN_445;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_24 <= _GEN_2748;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_25 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_25 <= _GEN_446;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_25 <= _GEN_2749;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_26 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_26 <= _GEN_447;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_26 <= _GEN_2750;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_27 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_27 <= _GEN_448;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_27 <= _GEN_2751;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_28 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_28 <= _GEN_449;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_28 <= _GEN_2752;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_29 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_29 <= _GEN_450;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_29 <= _GEN_2753;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_30 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_30 <= _GEN_451;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_30 <= _GEN_2754;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_31 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_31 <= _GEN_452;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_31 <= _GEN_2755;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_32 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_32 <= _GEN_453;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_32 <= _GEN_2756;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_33 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_33 <= _GEN_454;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_33 <= _GEN_2757;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_34 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_34 <= _GEN_455;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_34 <= _GEN_2758;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_35 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_35 <= _GEN_456;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_35 <= _GEN_2759;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_36 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_36 <= _GEN_457;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_36 <= _GEN_2760;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_37 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_37 <= _GEN_458;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_37 <= _GEN_2761;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_38 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_38 <= _GEN_459;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_38 <= _GEN_2762;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_39 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_39 <= _GEN_460;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_39 <= _GEN_2763;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_40 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_40 <= _GEN_461;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_40 <= _GEN_2764;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_41 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_41 <= _GEN_462;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_41 <= _GEN_2765;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_42 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_42 <= _GEN_463;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_42 <= _GEN_2766;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_43 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_43 <= _GEN_464;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_43 <= _GEN_2767;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_44 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_44 <= _GEN_465;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_44 <= _GEN_2768;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_45 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_45 <= _GEN_466;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_45 <= _GEN_2769;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_46 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_46 <= _GEN_467;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_46 <= _GEN_2770;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_47 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_47 <= _GEN_468;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_47 <= _GEN_2771;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_48 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_48 <= _GEN_469;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_48 <= _GEN_2772;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_49 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_49 <= _GEN_470;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_49 <= _GEN_2773;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_50 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_50 <= _GEN_471;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_50 <= _GEN_2774;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_51 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_51 <= _GEN_472;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_51 <= _GEN_2775;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_52 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_52 <= _GEN_473;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_52 <= _GEN_2776;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_53 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_53 <= _GEN_474;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_53 <= _GEN_2777;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_54 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_54 <= _GEN_475;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_54 <= _GEN_2778;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_55 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_55 <= _GEN_476;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_55 <= _GEN_2779;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_56 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_56 <= _GEN_477;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_56 <= _GEN_2780;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_57 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_57 <= _GEN_478;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_57 <= _GEN_2781;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_58 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_58 <= _GEN_479;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_58 <= _GEN_2782;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_59 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_59 <= _GEN_480;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_59 <= _GEN_2783;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_60 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_60 <= _GEN_481;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_60 <= _GEN_2784;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_61 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_61 <= _GEN_482;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_61 <= _GEN_2785;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_62 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_62 <= _GEN_483;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_62 <= _GEN_2786;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_63 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_63 <= _GEN_484;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_63 <= _GEN_2787;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_0 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_0 <= _GEN_485;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_0 <= _GEN_2788;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_1 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_1 <= _GEN_486;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_1 <= _GEN_2789;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_2 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_2 <= _GEN_487;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_2 <= _GEN_2790;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_3 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_3 <= _GEN_488;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_3 <= _GEN_2791;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_4 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_4 <= _GEN_489;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_4 <= _GEN_2792;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_5 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_5 <= _GEN_490;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_5 <= _GEN_2793;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_6 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_6 <= _GEN_491;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_6 <= _GEN_2794;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_7 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_7 <= _GEN_492;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_7 <= _GEN_2795;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_8 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_8 <= _GEN_493;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_8 <= _GEN_2796;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_9 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_9 <= _GEN_494;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_9 <= _GEN_2797;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_10 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_10 <= _GEN_495;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_10 <= _GEN_2798;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_11 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_11 <= _GEN_496;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_11 <= _GEN_2799;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_12 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_12 <= _GEN_497;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_12 <= _GEN_2800;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_13 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_13 <= _GEN_498;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_13 <= _GEN_2801;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_14 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_14 <= _GEN_499;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_14 <= _GEN_2802;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_15 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_15 <= _GEN_500;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_15 <= _GEN_2803;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_16 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_16 <= _GEN_501;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_16 <= _GEN_2804;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_17 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_17 <= _GEN_502;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_17 <= _GEN_2805;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_18 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_18 <= _GEN_503;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_18 <= _GEN_2806;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_19 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_19 <= _GEN_504;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_19 <= _GEN_2807;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_20 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_20 <= _GEN_505;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_20 <= _GEN_2808;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_21 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_21 <= _GEN_506;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_21 <= _GEN_2809;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_22 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_22 <= _GEN_507;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_22 <= _GEN_2810;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_23 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_23 <= _GEN_508;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_23 <= _GEN_2811;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_24 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_24 <= _GEN_509;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_24 <= _GEN_2812;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_25 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_25 <= _GEN_510;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_25 <= _GEN_2813;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_26 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_26 <= _GEN_511;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_26 <= _GEN_2814;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_27 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_27 <= _GEN_512;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_27 <= _GEN_2815;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_28 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_28 <= _GEN_513;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_28 <= _GEN_2816;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_29 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_29 <= _GEN_514;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_29 <= _GEN_2817;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_30 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_30 <= _GEN_515;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_30 <= _GEN_2818;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_31 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_31 <= _GEN_516;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_31 <= _GEN_2819;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_32 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_32 <= _GEN_517;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_32 <= _GEN_2820;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_33 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_33 <= _GEN_518;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_33 <= _GEN_2821;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_34 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_34 <= _GEN_519;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_34 <= _GEN_2822;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_35 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_35 <= _GEN_520;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_35 <= _GEN_2823;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_36 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_36 <= _GEN_521;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_36 <= _GEN_2824;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_37 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_37 <= _GEN_522;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_37 <= _GEN_2825;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_38 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_38 <= _GEN_523;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_38 <= _GEN_2826;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_39 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_39 <= _GEN_524;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_39 <= _GEN_2827;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_40 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_40 <= _GEN_525;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_40 <= _GEN_2828;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_41 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_41 <= _GEN_526;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_41 <= _GEN_2829;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_42 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_42 <= _GEN_527;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_42 <= _GEN_2830;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_43 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_43 <= _GEN_528;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_43 <= _GEN_2831;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_44 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_44 <= _GEN_529;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_44 <= _GEN_2832;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_45 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_45 <= _GEN_530;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_45 <= _GEN_2833;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_46 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_46 <= _GEN_531;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_46 <= _GEN_2834;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_47 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_47 <= _GEN_532;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_47 <= _GEN_2835;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_48 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_48 <= _GEN_533;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_48 <= _GEN_2836;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_49 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_49 <= _GEN_534;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_49 <= _GEN_2837;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_50 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_50 <= _GEN_535;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_50 <= _GEN_2838;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_51 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_51 <= _GEN_536;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_51 <= _GEN_2839;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_52 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_52 <= _GEN_537;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_52 <= _GEN_2840;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_53 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_53 <= _GEN_538;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_53 <= _GEN_2841;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_54 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_54 <= _GEN_539;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_54 <= _GEN_2842;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_55 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_55 <= _GEN_540;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_55 <= _GEN_2843;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_56 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_56 <= _GEN_541;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_56 <= _GEN_2844;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_57 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_57 <= _GEN_542;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_57 <= _GEN_2845;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_58 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_58 <= _GEN_543;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_58 <= _GEN_2846;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_59 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_59 <= _GEN_544;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_59 <= _GEN_2847;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_60 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_60 <= _GEN_545;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_60 <= _GEN_2848;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_61 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_61 <= _GEN_546;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_61 <= _GEN_2849;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_62 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_62 <= _GEN_547;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_62 <= _GEN_2850;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_63 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_63 <= _GEN_548;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_63 <= _GEN_2851;
      end
    end
    s2_hit_real_REG <= (hit_ready | _hit_ready_T) & io_in_resp_ready | invalid_ready; // @[Cache.scala 270:66]
    if (reset) begin // @[Cache.scala 209:25]
      s2_addr <= 32'h0; // @[Cache.scala 209:25]
    end else if (fi_ready) begin // @[Cache.scala 238:24]
      s2_addr <= io_in_req_bits_addr; // @[Cache.scala 240:14]
    end
    if (reset) begin // @[Cache.scala 231:27]
      s2_reg_hit <= 1'h0; // @[Cache.scala 231:27]
    end else if (!(fi_ready)) begin // @[Cache.scala 238:24]
      if (~fi_ready & REG) begin // @[Cache.scala 244:58]
        s2_reg_hit <= s2_hit; // @[Cache.scala 247:18]
      end
    end
    if (reset) begin // @[Cache.scala 213:25]
      s2_wen <= 1'h0; // @[Cache.scala 213:25]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      s2_wen <= _GEN_27;
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      s2_wen <= _GEN_27;
    end else if (_T_13) begin // @[Conditional.scala 39:67]
      s2_wen <= _GEN_27;
    end else begin
      s2_wen <= _GEN_2852;
    end
    if (reset) begin // @[Cache.scala 207:22]
      state <= 4'h8; // @[Cache.scala 207:22]
    end else if (fi_fire) begin // @[Cache.scala 411:18]
      state <= 4'h8; // @[Cache.scala 412:11]
    end else if (fi_ready) begin // @[Cache.scala 381:24]
      if (io_in_req_valid) begin // @[Cache.scala 382:17]
        state <= 4'h0;
      end else begin
        state <= 4'h8;
      end
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      state <= _GEN_983;
    end else begin
      state <= _GEN_3075;
    end
    if (reset) begin // @[ID.scala 18:20]
      fi_valid <= 1'h0; // @[ID.scala 18:20]
    end else if (dcache_fi_complete_0) begin // @[ID.scala 25:19]
      fi_valid <= 1'h0; // @[ID.scala 25:23]
    end else begin
      fi_valid <= _GEN_0;
    end
    if (reset) begin // @[Cache.scala 214:25]
      s2_wdata <= 64'h0; // @[Cache.scala 214:25]
    end else if (fi_ready) begin // @[Cache.scala 238:24]
      s2_wdata <= io_in_req_bits_wdata; // @[Cache.scala 242:14]
    end
    if (reset) begin // @[Cache.scala 215:25]
      s2_wmask <= 8'h0; // @[Cache.scala 215:25]
    end else if (fi_ready) begin // @[Cache.scala 238:24]
      s2_wmask <= io_in_req_bits_wmask; // @[Cache.scala 243:14]
    end
    if (reset) begin // @[Cache.scala 233:29]
      s2_reg_rdata <= 128'h0; // @[Cache.scala 233:29]
    end else if (!(fi_ready)) begin // @[Cache.scala 238:24]
      if (~fi_ready & REG) begin // @[Cache.scala 244:58]
        if (2'h3 == s2_way) begin // @[Cache.scala 249:18]
          s2_reg_rdata <= sram_out_3; // @[Cache.scala 249:18]
        end else begin
          s2_reg_rdata <= _GEN_6;
        end
      end
    end
    if (reset) begin // @[Cache.scala 234:29]
      s2_reg_dirty <= 1'h0; // @[Cache.scala 234:29]
    end else if (!(fi_ready)) begin // @[Cache.scala 238:24]
      if (~fi_ready & REG) begin // @[Cache.scala 244:58]
        if (2'h3 == replace_way) begin // @[Cache.scala 250:18]
          s2_reg_dirty <= dirty_out_3; // @[Cache.scala 250:18]
        end else begin
          s2_reg_dirty <= _GEN_10;
        end
      end
    end
    if (reset) begin // @[Cache.scala 235:29]
      s2_reg_tag_r <= 21'h0; // @[Cache.scala 235:29]
    end else if (!(fi_ready)) begin // @[Cache.scala 238:24]
      if (~fi_ready & REG) begin // @[Cache.scala 244:58]
        if (2'h3 == replace_way) begin // @[Cache.scala 251:18]
          s2_reg_tag_r <= tag_out_3; // @[Cache.scala 251:18]
        end else begin
          s2_reg_tag_r <= _GEN_14;
        end
      end
    end
    if (reset) begin // @[Cache.scala 236:29]
      s2_reg_dat_w <= 128'h0; // @[Cache.scala 236:29]
    end else if (!(fi_ready)) begin // @[Cache.scala 238:24]
      if (~fi_ready & REG) begin // @[Cache.scala 244:58]
        if (2'h3 == replace_way) begin // @[Cache.scala 252:18]
          s2_reg_dat_w <= sram_out_3; // @[Cache.scala 252:18]
        end else begin
          s2_reg_dat_w <= _GEN_18;
        end
      end
    end
    REG <= (hit_ready | _hit_ready_T) & io_in_resp_ready | invalid_ready; // @[Cache.scala 270:66]
    if (reset) begin // @[Cache.scala 258:23]
      wdata1 <= 64'h0; // @[Cache.scala 258:23]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (!(_T_11)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          wdata1 <= _GEN_988;
        end
      end
    end
    if (reset) begin // @[Cache.scala 259:23]
      wdata2 <= 64'h0; // @[Cache.scala 259:23]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (!(_T_11)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          wdata2 <= _GEN_989;
        end
      end
    end
    REG_1 <= (hit_ready | _hit_ready_T) & io_in_resp_ready | invalid_ready; // @[Cache.scala 270:66]
    REG_2 <= (hit_ready | _hit_ready_T) & io_in_resp_ready | invalid_ready; // @[Cache.scala 270:66]
    if (s2_offs) begin // @[Cache.scala 374:40]
      io_in_resp_bits_rdata_REG <= wdata2;
    end else begin
      io_in_resp_bits_rdata_REG <= wdata1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  plru0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  plru0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  plru0_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  plru0_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  plru0_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  plru0_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  plru0_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  plru0_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  plru0_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  plru0_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  plru0_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  plru0_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  plru0_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  plru0_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  plru0_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  plru0_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  plru0_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  plru0_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  plru0_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  plru0_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  plru0_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  plru0_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  plru0_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  plru0_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  plru0_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  plru0_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  plru0_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  plru0_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  plru0_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  plru0_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  plru0_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  plru0_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  plru0_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  plru0_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  plru0_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  plru0_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  plru0_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  plru0_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  plru0_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  plru0_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  plru0_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  plru0_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  plru0_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  plru0_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  plru0_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  plru0_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  plru0_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  plru0_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  plru0_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  plru0_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  plru0_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  plru0_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  plru0_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  plru0_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  plru0_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  plru0_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  plru0_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  plru0_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  plru0_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  plru0_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  plru0_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  plru0_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  plru0_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  plru0_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  plru1_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  plru1_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  plru1_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  plru1_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  plru1_4 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  plru1_5 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  plru1_6 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  plru1_7 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  plru1_8 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  plru1_9 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  plru1_10 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  plru1_11 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  plru1_12 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  plru1_13 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  plru1_14 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  plru1_15 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  plru1_16 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  plru1_17 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  plru1_18 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  plru1_19 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  plru1_20 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  plru1_21 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  plru1_22 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  plru1_23 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  plru1_24 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  plru1_25 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  plru1_26 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  plru1_27 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  plru1_28 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  plru1_29 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  plru1_30 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  plru1_31 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  plru1_32 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  plru1_33 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  plru1_34 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  plru1_35 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  plru1_36 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  plru1_37 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  plru1_38 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  plru1_39 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  plru1_40 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  plru1_41 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  plru1_42 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  plru1_43 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  plru1_44 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  plru1_45 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  plru1_46 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  plru1_47 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  plru1_48 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  plru1_49 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  plru1_50 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  plru1_51 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  plru1_52 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  plru1_53 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  plru1_54 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  plru1_55 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  plru1_56 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  plru1_57 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  plru1_58 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  plru1_59 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  plru1_60 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  plru1_61 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  plru1_62 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  plru1_63 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  plru2_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  plru2_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  plru2_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  plru2_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  plru2_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  plru2_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  plru2_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  plru2_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  plru2_8 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  plru2_9 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  plru2_10 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  plru2_11 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  plru2_12 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  plru2_13 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  plru2_14 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  plru2_15 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  plru2_16 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  plru2_17 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  plru2_18 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  plru2_19 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  plru2_20 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  plru2_21 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  plru2_22 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  plru2_23 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  plru2_24 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  plru2_25 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  plru2_26 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  plru2_27 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  plru2_28 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  plru2_29 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  plru2_30 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  plru2_31 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  plru2_32 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  plru2_33 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  plru2_34 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  plru2_35 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  plru2_36 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  plru2_37 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  plru2_38 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  plru2_39 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  plru2_40 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  plru2_41 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  plru2_42 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  plru2_43 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  plru2_44 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  plru2_45 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  plru2_46 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  plru2_47 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  plru2_48 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  plru2_49 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  plru2_50 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  plru2_51 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  plru2_52 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  plru2_53 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  plru2_54 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  plru2_55 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  plru2_56 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  plru2_57 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  plru2_58 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  plru2_59 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  plru2_60 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  plru2_61 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  plru2_62 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  plru2_63 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  s2_hit_real_REG = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  s2_addr = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  s2_reg_hit = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  s2_wen = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  state = _RAND_196[3:0];
  _RAND_197 = {1{`RANDOM}};
  fi_valid = _RAND_197[0:0];
  _RAND_198 = {2{`RANDOM}};
  s2_wdata = _RAND_198[63:0];
  _RAND_199 = {1{`RANDOM}};
  s2_wmask = _RAND_199[7:0];
  _RAND_200 = {4{`RANDOM}};
  s2_reg_rdata = _RAND_200[127:0];
  _RAND_201 = {1{`RANDOM}};
  s2_reg_dirty = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  s2_reg_tag_r = _RAND_202[20:0];
  _RAND_203 = {4{`RANDOM}};
  s2_reg_dat_w = _RAND_203[127:0];
  _RAND_204 = {1{`RANDOM}};
  REG = _RAND_204[0:0];
  _RAND_205 = {2{`RANDOM}};
  wdata1 = _RAND_205[63:0];
  _RAND_206 = {2{`RANDOM}};
  wdata2 = _RAND_206[63:0];
  _RAND_207 = {1{`RANDOM}};
  REG_1 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  REG_2 = _RAND_208[0:0];
  _RAND_209 = {2{`RANDOM}};
  io_in_resp_bits_rdata_REG = _RAND_209[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210340_Uncache(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input         io_in_req_bits_ren,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input  [1:0]  io_in_req_bits_size,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output        io_out_req_bits_ren,
  output [63:0] io_out_req_bits_wdata,
  output [7:0]  io_out_req_bits_wmask,
  output        io_out_req_bits_wen,
  output [1:0]  io_out_req_bits_size,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[Uncache.scala 18:22]
  reg [31:0] addr; // @[Uncache.scala 21:22]
  reg  ren; // @[Uncache.scala 22:22]
  reg [63:0] wdata; // @[Uncache.scala 23:22]
  reg [7:0] wmask; // @[Uncache.scala 24:22]
  reg  wen; // @[Uncache.scala 25:22]
  reg [1:0] size; // @[Uncache.scala 26:22]
  reg [63:0] rdata_1; // @[Uncache.scala 29:24]
  reg [63:0] rdata_2; // @[Uncache.scala 30:24]
  wire  req_split = size == 2'h3; // @[Uncache.scala 34:22]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_2 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_5 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _state_T = req_split ? 3'h3 : 3'h5; // @[Uncache.scala 59:21]
  wire [63:0] _GEN_10 = _T_5 ? io_out_resp_bits_rdata : rdata_1; // @[Uncache.scala 57:30 Uncache.scala 58:17 Uncache.scala 29:24]
  wire [2:0] _GEN_11 = _T_5 ? _state_T : state; // @[Uncache.scala 57:30 Uncache.scala 59:15 Uncache.scala 18:22]
  wire  _T_6 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_12 = _T_3 ? 3'h4 : state; // @[Uncache.scala 63:29 Uncache.scala 64:15 Uncache.scala 18:22]
  wire  _T_8 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire [63:0] _GEN_13 = _T_5 ? io_out_resp_bits_rdata : rdata_2; // @[Uncache.scala 68:30 Uncache.scala 69:17 Uncache.scala 30:24]
  wire [2:0] _GEN_14 = _T_5 ? 3'h5 : state; // @[Uncache.scala 68:30 Uncache.scala 70:15 Uncache.scala 18:22]
  wire  _T_10 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_11 = io_in_resp_ready & io_in_resp_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_15 = _T_11 ? 3'h0 : state; // @[Uncache.scala 74:29 Uncache.scala 75:15 Uncache.scala 18:22]
  wire [2:0] _GEN_16 = _T_10 ? _GEN_15 : state; // @[Conditional.scala 39:67 Uncache.scala 18:22]
  wire [63:0] _GEN_17 = _T_8 ? _GEN_13 : rdata_2; // @[Conditional.scala 39:67 Uncache.scala 30:24]
  wire [2:0] _GEN_18 = _T_8 ? _GEN_14 : _GEN_16; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_19 = _T_6 ? _GEN_12 : _GEN_18; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_20 = _T_6 ? rdata_2 : _GEN_17; // @[Conditional.scala 39:67 Uncache.scala 30:24]
  wire  _io_out_req_valid_T_1 = state == 3'h3; // @[Uncache.scala 81:55]
  wire [31:0] io_in_resp_bits_rdata_hi = rdata_2[31:0]; // @[Uncache.scala 91:53]
  wire [31:0] io_in_resp_bits_rdata_lo = rdata_1[31:0]; // @[Uncache.scala 91:68]
  wire [63:0] _io_in_resp_bits_rdata_T = {io_in_resp_bits_rdata_hi,io_in_resp_bits_rdata_lo}; // @[Cat.scala 30:58]
  wire [31:0] _io_out_req_bits_addr_T_3 = addr + 32'h4; // @[Uncache.scala 94:70]
  assign io_in_req_ready = state == 3'h0; // @[Uncache.scala 80:34]
  assign io_in_resp_valid = state == 3'h5; // @[Uncache.scala 90:34]
  assign io_in_resp_bits_rdata = req_split ? _io_in_resp_bits_rdata_T : rdata_1; // @[Uncache.scala 91:30]
  assign io_out_req_valid = state == 3'h1 | state == 3'h3; // @[Uncache.scala 81:46]
  assign io_out_req_bits_addr = req_split & _io_out_req_valid_T_1 ? _io_out_req_bits_addr_T_3 : addr; // @[Uncache.scala 94:30]
  assign io_out_req_bits_ren = ren; // @[Uncache.scala 84:24]
  assign io_out_req_bits_wdata = wdata; // @[Uncache.scala 95:24]
  assign io_out_req_bits_wmask = wmask; // @[Uncache.scala 96:24]
  assign io_out_req_bits_wen = wen; // @[Uncache.scala 86:24]
  assign io_out_req_bits_size = req_split ? 2'h2 : size; // @[Uncache.scala 97:30]
  assign io_out_resp_ready = state == 3'h2 | state == 3'h4; // @[Uncache.scala 89:47]
  always @(posedge clock) begin
    if (reset) begin // @[Uncache.scala 18:22]
      state <= 3'h0; // @[Uncache.scala 18:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        state <= 3'h1; // @[Uncache.scala 47:17]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Uncache.scala 52:29]
        state <= 3'h2; // @[Uncache.scala 53:15]
      end
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      state <= _GEN_11;
    end else begin
      state <= _GEN_19;
    end
    if (reset) begin // @[Uncache.scala 21:22]
      addr <= 32'h0; // @[Uncache.scala 21:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        addr <= io_in_req_bits_addr; // @[Uncache.scala 39:15]
      end
    end
    if (reset) begin // @[Uncache.scala 22:22]
      ren <= 1'h0; // @[Uncache.scala 22:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        ren <= io_in_req_bits_ren; // @[Uncache.scala 40:15]
      end
    end
    if (reset) begin // @[Uncache.scala 23:22]
      wdata <= 64'h0; // @[Uncache.scala 23:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        wdata <= io_in_req_bits_wdata; // @[Uncache.scala 41:15]
      end
    end
    if (reset) begin // @[Uncache.scala 24:22]
      wmask <= 8'h0; // @[Uncache.scala 24:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        wmask <= io_in_req_bits_wmask; // @[Uncache.scala 42:15]
      end
    end
    if (reset) begin // @[Uncache.scala 25:22]
      wen <= 1'h0; // @[Uncache.scala 25:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        wen <= io_in_req_bits_wen; // @[Uncache.scala 43:15]
      end
    end
    if (reset) begin // @[Uncache.scala 26:22]
      size <= 2'h0; // @[Uncache.scala 26:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        size <= io_in_req_bits_size; // @[Uncache.scala 44:15]
      end
    end
    if (reset) begin // @[Uncache.scala 29:24]
      rdata_1 <= 64'h0; // @[Uncache.scala 29:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        rdata_1 <= 64'h0; // @[Uncache.scala 45:17]
      end
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_4) begin // @[Conditional.scala 39:67]
        rdata_1 <= _GEN_10;
      end
    end
    if (reset) begin // @[Uncache.scala 30:24]
      rdata_2 <= 64'h0; // @[Uncache.scala 30:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        rdata_2 <= 64'h0; // @[Uncache.scala 46:17]
      end
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        rdata_2 <= _GEN_20;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  ren = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  wdata = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  wmask = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  wen = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  size = _RAND_6[1:0];
  _RAND_7 = {2{`RANDOM}};
  rdata_1 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  rdata_2 = _RAND_8[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210340_RRArbiter(
  input         clock,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_rdata,
  input         io_in_1_valid,
  input  [63:0] io_in_1_bits_rdata,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_rdata,
  output        io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _ctrl_validMask_grantMask_lastGrant_T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg  lastGrant; // @[Reg.scala 15:16]
  wire  grantMask_1 = 1'h1 > lastGrant; // @[Arbiter.scala 67:49]
  wire  validMask_1 = io_in_1_valid & grantMask_1; // @[Arbiter.scala 68:75]
  wire  _GEN_5 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:27 Arbiter.scala 77:36]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16 Arbiter.scala 41:16]
  assign io_out_bits_rdata = io_chosen ? io_in_1_bits_rdata : io_in_0_bits_rdata; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_chosen = validMask_1 | _GEN_5; // @[Arbiter.scala 79:25 Arbiter.scala 79:34]
  always @(posedge clock) begin
    if (_ctrl_validMask_grantMask_lastGrant_T) begin // @[Reg.scala 16:19]
      lastGrant <= io_chosen; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lastGrant = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210340_CacheBusCrossbar1to2(
  input         clock,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input         io_in_req_bits_ren,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input  [1:0]  io_in_req_bits_size,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_0_req_ready,
  output        io_out_0_req_valid,
  output [31:0] io_out_0_req_bits_addr,
  output        io_out_0_req_bits_ren,
  output [63:0] io_out_0_req_bits_wdata,
  output [7:0]  io_out_0_req_bits_wmask,
  output        io_out_0_req_bits_wen,
  output [1:0]  io_out_0_req_bits_size,
  output        io_out_0_resp_ready,
  input         io_out_0_resp_valid,
  input  [63:0] io_out_0_resp_bits_rdata,
  input         io_out_1_req_ready,
  output        io_out_1_req_valid,
  output [31:0] io_out_1_req_bits_addr,
  output        io_out_1_req_bits_ren,
  output [63:0] io_out_1_req_bits_wdata,
  output [7:0]  io_out_1_req_bits_wmask,
  output        io_out_1_req_bits_wen,
  output [1:0]  io_out_1_req_bits_size,
  output        io_out_1_resp_ready,
  input         io_out_1_resp_valid,
  input  [63:0] io_out_1_resp_bits_rdata,
  input         io_to_1
);
  wire  arbiter_clock; // @[Crossbar.scala 66:23]
  wire  arbiter_io_in_0_valid; // @[Crossbar.scala 66:23]
  wire [63:0] arbiter_io_in_0_bits_rdata; // @[Crossbar.scala 66:23]
  wire  arbiter_io_in_1_valid; // @[Crossbar.scala 66:23]
  wire [63:0] arbiter_io_in_1_bits_rdata; // @[Crossbar.scala 66:23]
  wire  arbiter_io_out_ready; // @[Crossbar.scala 66:23]
  wire  arbiter_io_out_valid; // @[Crossbar.scala 66:23]
  wire [63:0] arbiter_io_out_bits_rdata; // @[Crossbar.scala 66:23]
  wire  arbiter_io_chosen; // @[Crossbar.scala 66:23]
  ysyx_210340_RRArbiter arbiter ( // @[Crossbar.scala 66:23]
    .clock(arbiter_clock),
    .io_in_0_valid(arbiter_io_in_0_valid),
    .io_in_0_bits_rdata(arbiter_io_in_0_bits_rdata),
    .io_in_1_valid(arbiter_io_in_1_valid),
    .io_in_1_bits_rdata(arbiter_io_in_1_bits_rdata),
    .io_out_ready(arbiter_io_out_ready),
    .io_out_valid(arbiter_io_out_valid),
    .io_out_bits_rdata(arbiter_io_out_bits_rdata),
    .io_chosen(arbiter_io_chosen)
  );
  assign io_in_req_ready = io_to_1 ? io_out_1_req_ready : io_out_0_req_ready; // @[Crossbar.scala 64:25]
  assign io_in_resp_valid = arbiter_io_out_valid; // @[Crossbar.scala 75:13]
  assign io_in_resp_bits_rdata = arbiter_io_out_bits_rdata; // @[Crossbar.scala 74:12]
  assign io_out_0_req_valid = io_in_req_valid & ~io_to_1; // @[Crossbar.scala 62:42]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 60:22]
  assign io_out_0_req_bits_ren = io_in_req_bits_ren; // @[Crossbar.scala 60:22]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 60:22]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 60:22]
  assign io_out_0_req_bits_wen = io_in_req_bits_wen; // @[Crossbar.scala 60:22]
  assign io_out_0_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 60:22]
  assign io_out_0_resp_ready = ~arbiter_io_chosen; // @[Crossbar.scala 71:46]
  assign io_out_1_req_valid = io_in_req_valid & io_to_1; // @[Crossbar.scala 63:42]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 61:22]
  assign io_out_1_req_bits_ren = io_in_req_bits_ren; // @[Crossbar.scala 61:22]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 61:22]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 61:22]
  assign io_out_1_req_bits_wen = io_in_req_bits_wen; // @[Crossbar.scala 61:22]
  assign io_out_1_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 61:22]
  assign io_out_1_resp_ready = arbiter_io_chosen; // @[Crossbar.scala 72:46]
  assign arbiter_clock = clock;
  assign arbiter_io_in_0_valid = io_out_0_resp_valid; // @[Crossbar.scala 67:20]
  assign arbiter_io_in_0_bits_rdata = io_out_0_resp_bits_rdata; // @[Crossbar.scala 67:20]
  assign arbiter_io_in_1_valid = io_out_1_resp_valid; // @[Crossbar.scala 68:20]
  assign arbiter_io_in_1_bits_rdata = io_out_1_resp_bits_rdata; // @[Crossbar.scala 68:20]
  assign arbiter_io_out_ready = io_in_resp_ready; // @[Crossbar.scala 76:13]
endmodule
module ysyx_210340_CacheController(
  input         clock,
  input         reset,
  output [5:0]   io_sram0_addr,
  output         io_sram0_cen,
  output         io_sram0_wen,
  output [127:0] io_sram0_wdata,
  input  [127:0] io_sram0_rdata,
  output [5:0]   io_sram1_addr,
  output         io_sram1_cen,
  output         io_sram1_wen,
  output [127:0] io_sram1_wdata,
  input  [127:0] io_sram1_rdata,
  output [5:0]   io_sram2_addr,
  output         io_sram2_cen,
  output         io_sram2_wen,
  output [127:0] io_sram2_wdata,
  input  [127:0] io_sram2_rdata,
  output [5:0]   io_sram3_addr,
  output         io_sram3_cen,
  output         io_sram3_wen,
  output [127:0] io_sram3_wdata,
  input  [127:0] io_sram3_rdata,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_cache_req_ready,
  output        io_out_cache_req_valid,
  output [31:0] io_out_cache_req_bits_addr,
  output        io_out_cache_req_bits_aen,
  output        io_out_cache_req_bits_ren,
  output [63:0] io_out_cache_req_bits_wdata,
  output        io_out_cache_req_bits_wlast,
  output        io_out_cache_req_bits_wen,
  output        io_out_cache_resp_ready,
  input         io_out_cache_resp_valid,
  input  [63:0] io_out_cache_resp_bits_rdata,
  input         io_out_cache_resp_bits_rlast,
  input         io_out_uncache_req_ready,
  output        io_out_uncache_req_valid,
  output [31:0] io_out_uncache_req_bits_addr,
  output        io_out_uncache_req_bits_ren,
  output [63:0] io_out_uncache_req_bits_wdata,
  output [7:0]  io_out_uncache_req_bits_wmask,
  output        io_out_uncache_req_bits_wen,
  output [1:0]  io_out_uncache_req_bits_size,
  output        io_out_uncache_resp_ready,
  input         io_out_uncache_resp_valid,
  input  [63:0] io_out_uncache_resp_bits_rdata,
  input         fence_i,
  input         dcache_fi_complete
);

  wire [5:0] icache_io_sram0_addr; 
  wire  icache_io_sram0_cen; 
  wire  icache_io_sram0_wen; 
  wire [127:0] icache_io_sram0_wdata; 
  wire [127:0] icache_io_sram0_rdata; 
  wire [5:0] icache_io_sram1_addr; 
  wire  icache_io_sram1_cen; 
  wire  icache_io_sram1_wen; 
  wire [127:0] icache_io_sram1_wdata; 
  wire [127:0] icache_io_sram1_rdata; 
  wire [5:0] icache_io_sram2_addr; 
  wire  icache_io_sram2_cen; 
  wire  icache_io_sram2_wen; 
  wire [127:0] icache_io_sram2_wdata; 
  wire [127:0] icache_io_sram2_rdata; 
  wire [5:0] icache_io_sram3_addr; 
  wire  icache_io_sram3_cen; 
  wire  icache_io_sram3_wen; 
  wire [127:0] icache_io_sram3_wdata; 
  wire [127:0] icache_io_sram3_rdata; 

  wire  cache_clock; // @[CacheController.scala 14:21]
  wire  cache_reset; // @[CacheController.scala 14:21]
  wire  cache_io_in_req_ready; // @[CacheController.scala 14:21]
  wire  cache_io_in_req_valid; // @[CacheController.scala 14:21]
  wire [31:0] cache_io_in_req_bits_addr; // @[CacheController.scala 14:21]
  wire [63:0] cache_io_in_req_bits_wdata; // @[CacheController.scala 14:21]
  wire [7:0] cache_io_in_req_bits_wmask; // @[CacheController.scala 14:21]
  wire  cache_io_in_req_bits_wen; // @[CacheController.scala 14:21]
  wire  cache_io_in_resp_ready; // @[CacheController.scala 14:21]
  wire  cache_io_in_resp_valid; // @[CacheController.scala 14:21]
  wire [63:0] cache_io_in_resp_bits_rdata; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_ready; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_valid; // @[CacheController.scala 14:21]
  wire [31:0] cache_io_out_req_bits_addr; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_bits_aen; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_bits_ren; // @[CacheController.scala 14:21]
  wire [63:0] cache_io_out_req_bits_wdata; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_bits_wlast; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_bits_wen; // @[CacheController.scala 14:21]
  wire  cache_io_out_resp_ready; // @[CacheController.scala 14:21]
  wire  cache_io_out_resp_valid; // @[CacheController.scala 14:21]
  wire [63:0] cache_io_out_resp_bits_rdata; // @[CacheController.scala 14:21]
  wire  cache_io_out_resp_bits_rlast; // @[CacheController.scala 14:21]
  wire  cache_fence_i_0; // @[CacheController.scala 14:21]
  wire  cache_dcache_fi_complete_0; // @[CacheController.scala 14:21]
  wire  uncache_clock; // @[CacheController.scala 15:23]
  wire  uncache_reset; // @[CacheController.scala 15:23]
  wire  uncache_io_in_req_ready; // @[CacheController.scala 15:23]
  wire  uncache_io_in_req_valid; // @[CacheController.scala 15:23]
  wire [31:0] uncache_io_in_req_bits_addr; // @[CacheController.scala 15:23]
  wire  uncache_io_in_req_bits_ren; // @[CacheController.scala 15:23]
  wire [63:0] uncache_io_in_req_bits_wdata; // @[CacheController.scala 15:23]
  wire [7:0] uncache_io_in_req_bits_wmask; // @[CacheController.scala 15:23]
  wire  uncache_io_in_req_bits_wen; // @[CacheController.scala 15:23]
  wire [1:0] uncache_io_in_req_bits_size; // @[CacheController.scala 15:23]
  wire  uncache_io_in_resp_ready; // @[CacheController.scala 15:23]
  wire  uncache_io_in_resp_valid; // @[CacheController.scala 15:23]
  wire [63:0] uncache_io_in_resp_bits_rdata; // @[CacheController.scala 15:23]
  wire  uncache_io_out_req_ready; // @[CacheController.scala 15:23]
  wire  uncache_io_out_req_valid; // @[CacheController.scala 15:23]
  wire [31:0] uncache_io_out_req_bits_addr; // @[CacheController.scala 15:23]
  wire  uncache_io_out_req_bits_ren; // @[CacheController.scala 15:23]
  wire [63:0] uncache_io_out_req_bits_wdata; // @[CacheController.scala 15:23]
  wire [7:0] uncache_io_out_req_bits_wmask; // @[CacheController.scala 15:23]
  wire  uncache_io_out_req_bits_wen; // @[CacheController.scala 15:23]
  wire [1:0] uncache_io_out_req_bits_size; // @[CacheController.scala 15:23]
  wire  uncache_io_out_resp_ready; // @[CacheController.scala 15:23]
  wire  uncache_io_out_resp_valid; // @[CacheController.scala 15:23]
  wire [63:0] uncache_io_out_resp_bits_rdata; // @[CacheController.scala 15:23]
  wire  crossbar1to2_clock; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_req_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_req_valid; // @[CacheController.scala 17:28]
  wire [31:0] crossbar1to2_io_in_req_bits_addr; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_req_bits_ren; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_in_req_bits_wdata; // @[CacheController.scala 17:28]
  wire [7:0] crossbar1to2_io_in_req_bits_wmask; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_req_bits_wen; // @[CacheController.scala 17:28]
  wire [1:0] crossbar1to2_io_in_req_bits_size; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_resp_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_resp_valid; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_in_resp_bits_rdata; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_req_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_req_valid; // @[CacheController.scala 17:28]
  wire [31:0] crossbar1to2_io_out_0_req_bits_addr; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_req_bits_ren; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_out_0_req_bits_wdata; // @[CacheController.scala 17:28]
  wire [7:0] crossbar1to2_io_out_0_req_bits_wmask; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_req_bits_wen; // @[CacheController.scala 17:28]
  wire [1:0] crossbar1to2_io_out_0_req_bits_size; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_resp_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_resp_valid; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_out_0_resp_bits_rdata; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_req_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_req_valid; // @[CacheController.scala 17:28]
  wire [31:0] crossbar1to2_io_out_1_req_bits_addr; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_req_bits_ren; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_out_1_req_bits_wdata; // @[CacheController.scala 17:28]
  wire [7:0] crossbar1to2_io_out_1_req_bits_wmask; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_req_bits_wen; // @[CacheController.scala 17:28]
  wire [1:0] crossbar1to2_io_out_1_req_bits_size; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_resp_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_resp_valid; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_out_1_resp_bits_rdata; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_to_1; // @[CacheController.scala 17:28]
  ysyx_210340_Cache cache ( // @[CacheController.scala 14:21]
    .clock(cache_clock),
    .reset(cache_reset),
    .io_sram0_cen(icache_io_sram0_cen), 
    .io_sram0_wen(icache_io_sram0_wen), 
    .io_sram0_addr(icache_io_sram0_addr), 
    .io_sram0_wdata(icache_io_sram0_wdata), 
    .io_sram0_rdata(icache_io_sram0_rdata), 
    .io_sram1_cen(icache_io_sram1_cen), 
    .io_sram1_wen(icache_io_sram1_wen), 
    .io_sram1_addr(icache_io_sram1_addr), 
    .io_sram1_wdata(icache_io_sram1_wdata), 
    .io_sram1_rdata(icache_io_sram1_rdata),  
    .io_sram2_cen(icache_io_sram2_cen), 
    .io_sram2_wen(icache_io_sram2_wen), 
    .io_sram2_addr(icache_io_sram2_addr), 
    .io_sram2_wdata(icache_io_sram2_wdata), 
    .io_sram2_rdata(icache_io_sram2_rdata),   
    .io_sram3_cen(icache_io_sram3_cen), 
    .io_sram3_wen(icache_io_sram3_wen), 
    .io_sram3_addr(icache_io_sram3_addr), 
    .io_sram3_wdata(icache_io_sram3_wdata), 
    .io_sram3_rdata(icache_io_sram3_rdata),  
    .io_in_req_ready(cache_io_in_req_ready),
    .io_in_req_valid(cache_io_in_req_valid),
    .io_in_req_bits_addr(cache_io_in_req_bits_addr),
    .io_in_req_bits_wdata(cache_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(cache_io_in_req_bits_wmask),
    .io_in_req_bits_wen(cache_io_in_req_bits_wen),
    .io_in_resp_ready(cache_io_in_resp_ready),
    .io_in_resp_valid(cache_io_in_resp_valid),
    .io_in_resp_bits_rdata(cache_io_in_resp_bits_rdata),
    .io_out_req_ready(cache_io_out_req_ready),
    .io_out_req_valid(cache_io_out_req_valid),
    .io_out_req_bits_addr(cache_io_out_req_bits_addr),
    .io_out_req_bits_aen(cache_io_out_req_bits_aen),
    .io_out_req_bits_ren(cache_io_out_req_bits_ren),
    .io_out_req_bits_wdata(cache_io_out_req_bits_wdata),
    .io_out_req_bits_wlast(cache_io_out_req_bits_wlast),
    .io_out_req_bits_wen(cache_io_out_req_bits_wen),
    .io_out_resp_ready(cache_io_out_resp_ready),
    .io_out_resp_valid(cache_io_out_resp_valid),
    .io_out_resp_bits_rdata(cache_io_out_resp_bits_rdata),
    .io_out_resp_bits_rlast(cache_io_out_resp_bits_rlast),
    .fence_i_0(cache_fence_i_0),
    .dcache_fi_complete_0(cache_dcache_fi_complete_0)
  );

  assign io_sram0_addr = icache_io_sram0_addr; // @[cpu.scala 163:22]
  assign io_sram0_cen = icache_io_sram0_cen; // @[cpu.scala 163:22]
  assign io_sram0_wen = icache_io_sram0_wen; // @[cpu.scala 163:22]
  assign io_sram0_wdata = icache_io_sram0_wdata; // @[cpu.scala 163:22]
  assign io_sram1_addr = icache_io_sram1_addr; // @[cpu.scala 164:22]
  assign io_sram1_cen = icache_io_sram1_cen; // @[cpu.scala 164:22]
  assign io_sram1_wen = icache_io_sram1_wen; // @[cpu.scala 164:22]
  assign io_sram1_wdata = icache_io_sram1_wdata; // @[cpu.scala 164:22]
  assign io_sram2_addr = icache_io_sram2_addr; // @[cpu.scala 165:22]
  assign io_sram2_cen = icache_io_sram2_cen; // @[cpu.scala 165:22]
  assign io_sram2_wen = icache_io_sram2_wen; // @[cpu.scala 165:22]
  assign io_sram2_wdata = icache_io_sram2_wdata; // @[cpu.scala 165:22]
  assign io_sram3_addr = icache_io_sram3_addr; // @[cpu.scala 166:22]
  assign io_sram3_cen = icache_io_sram3_cen; // @[cpu.scala 166:22]
  assign io_sram3_wen = icache_io_sram3_wen; // @[cpu.scala 166:22]
  assign io_sram3_wdata = icache_io_sram3_wdata; // @[cpu.scala 166:22]

  assign icache_io_sram0_rdata = io_sram0_rdata;
  assign icache_io_sram1_rdata = io_sram1_rdata;
  assign icache_io_sram2_rdata = io_sram2_rdata;
  assign icache_io_sram3_rdata = io_sram3_rdata;

  ysyx_210340_Uncache uncache ( // @[CacheController.scala 15:23]
    .clock(uncache_clock),
    .reset(uncache_reset),
    .io_in_req_ready(uncache_io_in_req_ready),
    .io_in_req_valid(uncache_io_in_req_valid),
    .io_in_req_bits_addr(uncache_io_in_req_bits_addr),
    .io_in_req_bits_ren(uncache_io_in_req_bits_ren),
    .io_in_req_bits_wdata(uncache_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(uncache_io_in_req_bits_wmask),
    .io_in_req_bits_wen(uncache_io_in_req_bits_wen),
    .io_in_req_bits_size(uncache_io_in_req_bits_size),
    .io_in_resp_ready(uncache_io_in_resp_ready),
    .io_in_resp_valid(uncache_io_in_resp_valid),
    .io_in_resp_bits_rdata(uncache_io_in_resp_bits_rdata),
    .io_out_req_ready(uncache_io_out_req_ready),
    .io_out_req_valid(uncache_io_out_req_valid),
    .io_out_req_bits_addr(uncache_io_out_req_bits_addr),
    .io_out_req_bits_ren(uncache_io_out_req_bits_ren),
    .io_out_req_bits_wdata(uncache_io_out_req_bits_wdata),
    .io_out_req_bits_wmask(uncache_io_out_req_bits_wmask),
    .io_out_req_bits_wen(uncache_io_out_req_bits_wen),
    .io_out_req_bits_size(uncache_io_out_req_bits_size),
    .io_out_resp_ready(uncache_io_out_resp_ready),
    .io_out_resp_valid(uncache_io_out_resp_valid),
    .io_out_resp_bits_rdata(uncache_io_out_resp_bits_rdata)
  );
  ysyx_210340_CacheBusCrossbar1to2 crossbar1to2 ( // @[CacheController.scala 17:28]
    .clock(crossbar1to2_clock),
    .io_in_req_ready(crossbar1to2_io_in_req_ready),
    .io_in_req_valid(crossbar1to2_io_in_req_valid),
    .io_in_req_bits_addr(crossbar1to2_io_in_req_bits_addr),
    .io_in_req_bits_ren(crossbar1to2_io_in_req_bits_ren),
    .io_in_req_bits_wdata(crossbar1to2_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(crossbar1to2_io_in_req_bits_wmask),
    .io_in_req_bits_wen(crossbar1to2_io_in_req_bits_wen),
    .io_in_req_bits_size(crossbar1to2_io_in_req_bits_size),
    .io_in_resp_ready(crossbar1to2_io_in_resp_ready),
    .io_in_resp_valid(crossbar1to2_io_in_resp_valid),
    .io_in_resp_bits_rdata(crossbar1to2_io_in_resp_bits_rdata),
    .io_out_0_req_ready(crossbar1to2_io_out_0_req_ready),
    .io_out_0_req_valid(crossbar1to2_io_out_0_req_valid),
    .io_out_0_req_bits_addr(crossbar1to2_io_out_0_req_bits_addr),
    .io_out_0_req_bits_ren(crossbar1to2_io_out_0_req_bits_ren),
    .io_out_0_req_bits_wdata(crossbar1to2_io_out_0_req_bits_wdata),
    .io_out_0_req_bits_wmask(crossbar1to2_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wen(crossbar1to2_io_out_0_req_bits_wen),
    .io_out_0_req_bits_size(crossbar1to2_io_out_0_req_bits_size),
    .io_out_0_resp_ready(crossbar1to2_io_out_0_resp_ready),
    .io_out_0_resp_valid(crossbar1to2_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(crossbar1to2_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(crossbar1to2_io_out_1_req_ready),
    .io_out_1_req_valid(crossbar1to2_io_out_1_req_valid),
    .io_out_1_req_bits_addr(crossbar1to2_io_out_1_req_bits_addr),
    .io_out_1_req_bits_ren(crossbar1to2_io_out_1_req_bits_ren),
    .io_out_1_req_bits_wdata(crossbar1to2_io_out_1_req_bits_wdata),
    .io_out_1_req_bits_wmask(crossbar1to2_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wen(crossbar1to2_io_out_1_req_bits_wen),
    .io_out_1_req_bits_size(crossbar1to2_io_out_1_req_bits_size),
    .io_out_1_resp_ready(crossbar1to2_io_out_1_resp_ready),
    .io_out_1_resp_valid(crossbar1to2_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(crossbar1to2_io_out_1_resp_bits_rdata),
    .io_to_1(crossbar1to2_io_to_1)
  );
  assign io_in_req_ready = crossbar1to2_io_in_req_ready; // @[CacheController.scala 19:22]
  assign io_in_resp_valid = crossbar1to2_io_in_resp_valid; // @[CacheController.scala 19:22]
  assign io_in_resp_bits_rdata = crossbar1to2_io_in_resp_bits_rdata; // @[CacheController.scala 19:22]
  assign io_out_cache_req_valid = cache_io_out_req_valid; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_addr = cache_io_out_req_bits_addr; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_aen = cache_io_out_req_bits_aen; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_ren = cache_io_out_req_bits_ren; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_wdata = cache_io_out_req_bits_wdata; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_wlast = cache_io_out_req_bits_wlast; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_wen = cache_io_out_req_bits_wen; // @[CacheController.scala 23:16]
  assign io_out_cache_resp_ready = cache_io_out_resp_ready; // @[CacheController.scala 23:16]
  assign io_out_uncache_req_valid = uncache_io_out_req_valid; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_addr = uncache_io_out_req_bits_addr; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_ren = uncache_io_out_req_bits_ren; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_wdata = uncache_io_out_req_bits_wdata; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_wmask = uncache_io_out_req_bits_wmask; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_wen = uncache_io_out_req_bits_wen; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_size = uncache_io_out_req_bits_size; // @[CacheController.scala 24:18]
  assign io_out_uncache_resp_ready = uncache_io_out_resp_ready; // @[CacheController.scala 24:18]
  assign cache_clock = clock;
  assign cache_reset = reset;
  assign cache_io_in_req_valid = crossbar1to2_io_out_0_req_valid; // @[CacheController.scala 20:26]
  assign cache_io_in_req_bits_addr = crossbar1to2_io_out_0_req_bits_addr; // @[CacheController.scala 20:26]
  assign cache_io_in_req_bits_wdata = crossbar1to2_io_out_0_req_bits_wdata; // @[CacheController.scala 20:26]
  assign cache_io_in_req_bits_wmask = crossbar1to2_io_out_0_req_bits_wmask; // @[CacheController.scala 20:26]
  assign cache_io_in_req_bits_wen = crossbar1to2_io_out_0_req_bits_wen; // @[CacheController.scala 20:26]
  assign cache_io_in_resp_ready = crossbar1to2_io_out_0_resp_ready; // @[CacheController.scala 20:26]
  assign cache_io_out_req_ready = io_out_cache_req_ready; // @[CacheController.scala 23:16]
  assign cache_io_out_resp_valid = io_out_cache_resp_valid; // @[CacheController.scala 23:16]
  assign cache_io_out_resp_bits_rdata = io_out_cache_resp_bits_rdata; // @[CacheController.scala 23:16]
  assign cache_io_out_resp_bits_rlast = io_out_cache_resp_bits_rlast; // @[CacheController.scala 23:16]
  assign cache_fence_i_0 = fence_i;
  assign cache_dcache_fi_complete_0 = dcache_fi_complete;
  assign uncache_clock = clock;
  assign uncache_reset = reset;
  assign uncache_io_in_req_valid = crossbar1to2_io_out_1_req_valid; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_addr = crossbar1to2_io_out_1_req_bits_addr; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_ren = crossbar1to2_io_out_1_req_bits_ren; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_wdata = crossbar1to2_io_out_1_req_bits_wdata; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_wmask = crossbar1to2_io_out_1_req_bits_wmask; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_wen = crossbar1to2_io_out_1_req_bits_wen; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_size = crossbar1to2_io_out_1_req_bits_size; // @[CacheController.scala 21:26]
  assign uncache_io_in_resp_ready = crossbar1to2_io_out_1_resp_ready; // @[CacheController.scala 21:26]
  assign uncache_io_out_req_ready = io_out_uncache_req_ready; // @[CacheController.scala 24:18]
  assign uncache_io_out_resp_valid = io_out_uncache_resp_valid; // @[CacheController.scala 24:18]
  assign uncache_io_out_resp_bits_rdata = io_out_uncache_resp_bits_rdata; // @[CacheController.scala 24:18]
  assign crossbar1to2_clock = clock;
  assign crossbar1to2_io_in_req_valid = io_in_req_valid; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_addr = io_in_req_bits_addr; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_ren = 1'h1; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_wdata = 64'h0; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_wmask = 8'h0; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_wen = 1'h0; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_size = 2'h3; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_resp_ready = io_in_resp_ready; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_out_0_req_ready = cache_io_in_req_ready; // @[CacheController.scala 20:26]
  assign crossbar1to2_io_out_0_resp_valid = cache_io_in_resp_valid; // @[CacheController.scala 20:26]
  assign crossbar1to2_io_out_0_resp_bits_rdata = cache_io_in_resp_bits_rdata; // @[CacheController.scala 20:26]
  assign crossbar1to2_io_out_1_req_ready = uncache_io_in_req_ready; // @[CacheController.scala 21:26]
  assign crossbar1to2_io_out_1_resp_valid = uncache_io_in_resp_valid; // @[CacheController.scala 21:26]
  assign crossbar1to2_io_out_1_resp_bits_rdata = uncache_io_in_resp_bits_rdata; // @[CacheController.scala 21:26]
  assign crossbar1to2_io_to_1 = ~io_in_req_bits_addr[31]; // @[CacheController.scala 13:45]
endmodule
module ysyx_210340_PipelineReg(
  input         clock,
  input         reset,
  input  [31:0] io_in_pc,
  input  [31:0] io_in_inst,
  input         io_in_imem_hs,
  output [31:0] io_out_pc,
  output [31:0] io_out_inst,
  output        io_out_imem_hs,
  input         io_flush,
  input         io_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_pc; // @[PipelineReg.scala 60:20]
  reg [31:0] reg_inst; // @[PipelineReg.scala 60:20]
  reg  reg_imem_hs; // @[PipelineReg.scala 60:20]
  assign io_out_pc = reg_pc; // @[PipelineReg.scala 68:10]
  assign io_out_inst = reg_inst; // @[PipelineReg.scala 68:10]
  assign io_out_imem_hs = reg_imem_hs; // @[PipelineReg.scala 68:10]
  always @(posedge clock) begin
    if (reset) begin // @[PipelineReg.scala 60:20]
      reg_pc <= 32'h0; // @[PipelineReg.scala 60:20]
    end else if (io_flush) begin // @[PipelineReg.scala 62:19]
      reg_pc <= 32'h0; // @[PipelineReg.scala 15:17]
    end else if (~io_stall) begin // @[PipelineReg.scala 64:27]
      reg_pc <= io_in_pc; // @[PipelineReg.scala 65:9]
    end
    if (reset) begin // @[PipelineReg.scala 60:20]
      reg_inst <= 32'h0; // @[PipelineReg.scala 60:20]
    end else if (io_flush) begin // @[PipelineReg.scala 62:19]
      reg_inst <= 32'h0; // @[PipelineReg.scala 16:17]
    end else if (~io_stall) begin // @[PipelineReg.scala 64:27]
      reg_inst <= io_in_inst; // @[PipelineReg.scala 65:9]
    end
    if (reset) begin // @[PipelineReg.scala 60:20]
      reg_imem_hs <= 1'h0; // @[PipelineReg.scala 60:20]
    end else if (io_flush) begin // @[PipelineReg.scala 62:19]
      reg_imem_hs <= 1'h0; // @[PipelineReg.scala 17:17]
    end else if (~io_stall) begin // @[PipelineReg.scala 64:27]
      reg_imem_hs <= io_in_imem_hs; // @[PipelineReg.scala 65:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_inst = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_imem_hs = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210340_Decode(
  input  [31:0] io_inst,
  output [4:0]  io_rs1_addr,
  output [1:0]  io_rs1_type,
  output [4:0]  io_rs2_addr,
  output [1:0]  io_rs2_type,
  output [4:0]  io_rd_addr,
  output        io_rd_en,
  output [5:0]  io_op_type,
  output [2:0]  io_fuType,
  output [63:0] io_imm,
  output [63:0] io_csr_imm
);
  wire [31:0] _T = io_inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _T_1 = 32'h13 == _T; // @[Lookup.scala 31:38]
  wire [31:0] _T_2 = io_inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _T_3 = 32'h1013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_5 = 32'h2013 == _T; // @[Lookup.scala 31:38]
  wire  _T_7 = 32'h3013 == _T; // @[Lookup.scala 31:38]
  wire  _T_9 = 32'h4013 == _T; // @[Lookup.scala 31:38]
  wire  _T_11 = 32'h5013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_13 = 32'h7013 == _T; // @[Lookup.scala 31:38]
  wire  _T_15 = 32'h40005013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_17 = 32'h6013 == _T; // @[Lookup.scala 31:38]
  wire [31:0] _T_18 = io_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _T_19 = 32'h33 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_21 = 32'h1033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_23 = 32'h2033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_25 = 32'h3033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_27 = 32'h4033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_29 = 32'h5033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_31 = 32'h6033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_33 = 32'h7033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_35 = 32'h40000033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_37 = 32'h40005033 == _T_18; // @[Lookup.scala 31:38]
  wire [31:0] _T_38 = io_inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _T_39 = 32'h17 == _T_38; // @[Lookup.scala 31:38]
  wire  _T_41 = 32'h37 == _T_38; // @[Lookup.scala 31:38]
  wire  _T_43 = 32'h1b == _T; // @[Lookup.scala 31:38]
  wire  _T_45 = 32'h101b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_47 = 32'h501b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_49 = 32'h4000501b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_51 = 32'h103b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_53 = 32'h503b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_55 = 32'h4000503b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_57 = 32'h3b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_59 = 32'h4000003b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_61 = 32'h6f == _T_38; // @[Lookup.scala 31:38]
  wire  _T_63 = 32'h67 == _T; // @[Lookup.scala 31:38]
  wire  _T_65 = 32'h63 == _T; // @[Lookup.scala 31:38]
  wire  _T_67 = 32'h1063 == _T; // @[Lookup.scala 31:38]
  wire  _T_69 = 32'h4063 == _T; // @[Lookup.scala 31:38]
  wire  _T_71 = 32'h5063 == _T; // @[Lookup.scala 31:38]
  wire  _T_73 = 32'h6063 == _T; // @[Lookup.scala 31:38]
  wire  _T_75 = 32'h7063 == _T; // @[Lookup.scala 31:38]
  wire  _T_77 = 32'h3 == _T; // @[Lookup.scala 31:38]
  wire  _T_79 = 32'h1003 == _T; // @[Lookup.scala 31:38]
  wire  _T_81 = 32'h2003 == _T; // @[Lookup.scala 31:38]
  wire  _T_83 = 32'h3003 == _T; // @[Lookup.scala 31:38]
  wire  _T_85 = 32'h4003 == _T; // @[Lookup.scala 31:38]
  wire  _T_87 = 32'h5003 == _T; // @[Lookup.scala 31:38]
  wire  _T_89 = 32'h6003 == _T; // @[Lookup.scala 31:38]
  wire  _T_91 = 32'h23 == _T; // @[Lookup.scala 31:38]
  wire  _T_93 = 32'h1023 == _T; // @[Lookup.scala 31:38]
  wire  _T_95 = 32'h2023 == _T; // @[Lookup.scala 31:38]
  wire  _T_97 = 32'h3023 == _T; // @[Lookup.scala 31:38]
  wire  _T_99 = 32'h1073 == _T; // @[Lookup.scala 31:38]
  wire  _T_101 = 32'h2073 == _T; // @[Lookup.scala 31:38]
  wire  _T_103 = 32'h3073 == _T; // @[Lookup.scala 31:38]
  wire  _T_105 = 32'h5073 == _T; // @[Lookup.scala 31:38]
  wire  _T_107 = 32'h6073 == _T; // @[Lookup.scala 31:38]
  wire  _T_109 = 32'h7073 == _T; // @[Lookup.scala 31:38]
  wire  _T_111 = 32'h73 == io_inst; // @[Lookup.scala 31:38]
  wire  _T_113 = 32'h30200073 == io_inst; // @[Lookup.scala 31:38]
  wire  _T_115 = 32'h13 == io_inst; // @[Lookup.scala 31:38]
  wire  _T_117 = 32'h100f == io_inst; // @[Lookup.scala 31:38]
  wire [2:0] _T_119 = _T_115 ? 3'h4 : {{2'd0}, _T_117}; // @[Lookup.scala 33:37]
  wire [2:0] _T_120 = _T_113 ? 3'h4 : _T_119; // @[Lookup.scala 33:37]
  wire [2:0] _T_121 = _T_111 ? 3'h4 : _T_120; // @[Lookup.scala 33:37]
  wire [2:0] _T_122 = _T_109 ? 3'h4 : _T_121; // @[Lookup.scala 33:37]
  wire [2:0] _T_123 = _T_107 ? 3'h4 : _T_122; // @[Lookup.scala 33:37]
  wire [2:0] _T_124 = _T_105 ? 3'h4 : _T_123; // @[Lookup.scala 33:37]
  wire [2:0] _T_125 = _T_103 ? 3'h4 : _T_124; // @[Lookup.scala 33:37]
  wire [2:0] _T_126 = _T_101 ? 3'h4 : _T_125; // @[Lookup.scala 33:37]
  wire [2:0] _T_127 = _T_99 ? 3'h4 : _T_126; // @[Lookup.scala 33:37]
  wire [2:0] _T_128 = _T_97 ? 3'h2 : _T_127; // @[Lookup.scala 33:37]
  wire [2:0] _T_129 = _T_95 ? 3'h2 : _T_128; // @[Lookup.scala 33:37]
  wire [2:0] _T_130 = _T_93 ? 3'h2 : _T_129; // @[Lookup.scala 33:37]
  wire [2:0] _T_131 = _T_91 ? 3'h2 : _T_130; // @[Lookup.scala 33:37]
  wire [2:0] _T_132 = _T_89 ? 3'h4 : _T_131; // @[Lookup.scala 33:37]
  wire [2:0] _T_133 = _T_87 ? 3'h4 : _T_132; // @[Lookup.scala 33:37]
  wire [2:0] _T_134 = _T_85 ? 3'h4 : _T_133; // @[Lookup.scala 33:37]
  wire [2:0] _T_135 = _T_83 ? 3'h4 : _T_134; // @[Lookup.scala 33:37]
  wire [2:0] _T_136 = _T_81 ? 3'h4 : _T_135; // @[Lookup.scala 33:37]
  wire [2:0] _T_137 = _T_79 ? 3'h4 : _T_136; // @[Lookup.scala 33:37]
  wire [2:0] _T_138 = _T_77 ? 3'h4 : _T_137; // @[Lookup.scala 33:37]
  wire [2:0] _T_139 = _T_75 ? 3'h1 : _T_138; // @[Lookup.scala 33:37]
  wire [2:0] _T_140 = _T_73 ? 3'h1 : _T_139; // @[Lookup.scala 33:37]
  wire [2:0] _T_141 = _T_71 ? 3'h1 : _T_140; // @[Lookup.scala 33:37]
  wire [2:0] _T_142 = _T_69 ? 3'h1 : _T_141; // @[Lookup.scala 33:37]
  wire [2:0] _T_143 = _T_67 ? 3'h1 : _T_142; // @[Lookup.scala 33:37]
  wire [2:0] _T_144 = _T_65 ? 3'h1 : _T_143; // @[Lookup.scala 33:37]
  wire [2:0] _T_145 = _T_63 ? 3'h4 : _T_144; // @[Lookup.scala 33:37]
  wire [2:0] _T_146 = _T_61 ? 3'h7 : _T_145; // @[Lookup.scala 33:37]
  wire [2:0] _T_147 = _T_59 ? 3'h5 : _T_146; // @[Lookup.scala 33:37]
  wire [2:0] _T_148 = _T_57 ? 3'h5 : _T_147; // @[Lookup.scala 33:37]
  wire [2:0] _T_149 = _T_55 ? 3'h5 : _T_148; // @[Lookup.scala 33:37]
  wire [2:0] _T_150 = _T_53 ? 3'h5 : _T_149; // @[Lookup.scala 33:37]
  wire [2:0] _T_151 = _T_51 ? 3'h5 : _T_150; // @[Lookup.scala 33:37]
  wire [2:0] _T_152 = _T_49 ? 3'h4 : _T_151; // @[Lookup.scala 33:37]
  wire [2:0] _T_153 = _T_47 ? 3'h4 : _T_152; // @[Lookup.scala 33:37]
  wire [2:0] _T_154 = _T_45 ? 3'h4 : _T_153; // @[Lookup.scala 33:37]
  wire [2:0] _T_155 = _T_43 ? 3'h4 : _T_154; // @[Lookup.scala 33:37]
  wire [2:0] _T_156 = _T_41 ? 3'h6 : _T_155; // @[Lookup.scala 33:37]
  wire [2:0] _T_157 = _T_39 ? 3'h6 : _T_156; // @[Lookup.scala 33:37]
  wire [2:0] _T_158 = _T_37 ? 3'h5 : _T_157; // @[Lookup.scala 33:37]
  wire [2:0] _T_159 = _T_35 ? 3'h5 : _T_158; // @[Lookup.scala 33:37]
  wire [2:0] _T_160 = _T_33 ? 3'h5 : _T_159; // @[Lookup.scala 33:37]
  wire [2:0] _T_161 = _T_31 ? 3'h5 : _T_160; // @[Lookup.scala 33:37]
  wire [2:0] _T_162 = _T_29 ? 3'h5 : _T_161; // @[Lookup.scala 33:37]
  wire [2:0] _T_163 = _T_27 ? 3'h5 : _T_162; // @[Lookup.scala 33:37]
  wire [2:0] _T_164 = _T_25 ? 3'h5 : _T_163; // @[Lookup.scala 33:37]
  wire [2:0] _T_165 = _T_23 ? 3'h5 : _T_164; // @[Lookup.scala 33:37]
  wire [2:0] _T_166 = _T_21 ? 3'h5 : _T_165; // @[Lookup.scala 33:37]
  wire [2:0] _T_167 = _T_19 ? 3'h5 : _T_166; // @[Lookup.scala 33:37]
  wire [2:0] _T_168 = _T_17 ? 3'h4 : _T_167; // @[Lookup.scala 33:37]
  wire [2:0] _T_169 = _T_15 ? 3'h4 : _T_168; // @[Lookup.scala 33:37]
  wire [2:0] _T_170 = _T_13 ? 3'h4 : _T_169; // @[Lookup.scala 33:37]
  wire [2:0] _T_171 = _T_11 ? 3'h4 : _T_170; // @[Lookup.scala 33:37]
  wire [2:0] _T_172 = _T_9 ? 3'h4 : _T_171; // @[Lookup.scala 33:37]
  wire [2:0] _T_173 = _T_7 ? 3'h4 : _T_172; // @[Lookup.scala 33:37]
  wire [2:0] _T_174 = _T_5 ? 3'h4 : _T_173; // @[Lookup.scala 33:37]
  wire [2:0] _T_175 = _T_3 ? 3'h4 : _T_174; // @[Lookup.scala 33:37]
  wire [2:0] instrType = _T_1 ? 3'h4 : _T_175; // @[Lookup.scala 33:37]
  wire [2:0] _T_176 = _T_117 ? 3'h4 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_177 = _T_115 ? 3'h0 : _T_176; // @[Lookup.scala 33:37]
  wire [2:0] _T_178 = _T_113 ? 3'h3 : _T_177; // @[Lookup.scala 33:37]
  wire [2:0] _T_179 = _T_111 ? 3'h3 : _T_178; // @[Lookup.scala 33:37]
  wire [2:0] _T_180 = _T_109 ? 3'h3 : _T_179; // @[Lookup.scala 33:37]
  wire [2:0] _T_181 = _T_107 ? 3'h3 : _T_180; // @[Lookup.scala 33:37]
  wire [2:0] _T_182 = _T_105 ? 3'h3 : _T_181; // @[Lookup.scala 33:37]
  wire [2:0] _T_183 = _T_103 ? 3'h3 : _T_182; // @[Lookup.scala 33:37]
  wire [2:0] _T_184 = _T_101 ? 3'h3 : _T_183; // @[Lookup.scala 33:37]
  wire [2:0] _T_185 = _T_99 ? 3'h3 : _T_184; // @[Lookup.scala 33:37]
  wire [2:0] _T_186 = _T_97 ? 3'h2 : _T_185; // @[Lookup.scala 33:37]
  wire [2:0] _T_187 = _T_95 ? 3'h2 : _T_186; // @[Lookup.scala 33:37]
  wire [2:0] _T_188 = _T_93 ? 3'h2 : _T_187; // @[Lookup.scala 33:37]
  wire [2:0] _T_189 = _T_91 ? 3'h2 : _T_188; // @[Lookup.scala 33:37]
  wire [2:0] _T_190 = _T_89 ? 3'h2 : _T_189; // @[Lookup.scala 33:37]
  wire [2:0] _T_191 = _T_87 ? 3'h2 : _T_190; // @[Lookup.scala 33:37]
  wire [2:0] _T_192 = _T_85 ? 3'h2 : _T_191; // @[Lookup.scala 33:37]
  wire [2:0] _T_193 = _T_83 ? 3'h2 : _T_192; // @[Lookup.scala 33:37]
  wire [2:0] _T_194 = _T_81 ? 3'h2 : _T_193; // @[Lookup.scala 33:37]
  wire [2:0] _T_195 = _T_79 ? 3'h2 : _T_194; // @[Lookup.scala 33:37]
  wire [2:0] _T_196 = _T_77 ? 3'h2 : _T_195; // @[Lookup.scala 33:37]
  wire [2:0] _T_197 = _T_75 ? 3'h1 : _T_196; // @[Lookup.scala 33:37]
  wire [2:0] _T_198 = _T_73 ? 3'h1 : _T_197; // @[Lookup.scala 33:37]
  wire [2:0] _T_199 = _T_71 ? 3'h1 : _T_198; // @[Lookup.scala 33:37]
  wire [2:0] _T_200 = _T_69 ? 3'h1 : _T_199; // @[Lookup.scala 33:37]
  wire [2:0] _T_201 = _T_67 ? 3'h1 : _T_200; // @[Lookup.scala 33:37]
  wire [2:0] _T_202 = _T_65 ? 3'h1 : _T_201; // @[Lookup.scala 33:37]
  wire [2:0] _T_203 = _T_63 ? 3'h1 : _T_202; // @[Lookup.scala 33:37]
  wire [2:0] _T_204 = _T_61 ? 3'h1 : _T_203; // @[Lookup.scala 33:37]
  wire [2:0] _T_205 = _T_59 ? 3'h0 : _T_204; // @[Lookup.scala 33:37]
  wire [2:0] _T_206 = _T_57 ? 3'h0 : _T_205; // @[Lookup.scala 33:37]
  wire [2:0] _T_207 = _T_55 ? 3'h0 : _T_206; // @[Lookup.scala 33:37]
  wire [2:0] _T_208 = _T_53 ? 3'h0 : _T_207; // @[Lookup.scala 33:37]
  wire [2:0] _T_209 = _T_51 ? 3'h0 : _T_208; // @[Lookup.scala 33:37]
  wire [2:0] _T_210 = _T_49 ? 3'h0 : _T_209; // @[Lookup.scala 33:37]
  wire [2:0] _T_211 = _T_47 ? 3'h0 : _T_210; // @[Lookup.scala 33:37]
  wire [2:0] _T_212 = _T_45 ? 3'h0 : _T_211; // @[Lookup.scala 33:37]
  wire [2:0] _T_213 = _T_43 ? 3'h0 : _T_212; // @[Lookup.scala 33:37]
  wire [2:0] _T_214 = _T_41 ? 3'h0 : _T_213; // @[Lookup.scala 33:37]
  wire [2:0] _T_215 = _T_39 ? 3'h0 : _T_214; // @[Lookup.scala 33:37]
  wire [2:0] _T_216 = _T_37 ? 3'h0 : _T_215; // @[Lookup.scala 33:37]
  wire [2:0] _T_217 = _T_35 ? 3'h0 : _T_216; // @[Lookup.scala 33:37]
  wire [2:0] _T_218 = _T_33 ? 3'h0 : _T_217; // @[Lookup.scala 33:37]
  wire [2:0] _T_219 = _T_31 ? 3'h0 : _T_218; // @[Lookup.scala 33:37]
  wire [2:0] _T_220 = _T_29 ? 3'h0 : _T_219; // @[Lookup.scala 33:37]
  wire [2:0] _T_221 = _T_27 ? 3'h0 : _T_220; // @[Lookup.scala 33:37]
  wire [2:0] _T_222 = _T_25 ? 3'h0 : _T_221; // @[Lookup.scala 33:37]
  wire [2:0] _T_223 = _T_23 ? 3'h0 : _T_222; // @[Lookup.scala 33:37]
  wire [2:0] _T_224 = _T_21 ? 3'h0 : _T_223; // @[Lookup.scala 33:37]
  wire [2:0] _T_225 = _T_19 ? 3'h0 : _T_224; // @[Lookup.scala 33:37]
  wire [2:0] _T_226 = _T_17 ? 3'h0 : _T_225; // @[Lookup.scala 33:37]
  wire [2:0] _T_227 = _T_15 ? 3'h0 : _T_226; // @[Lookup.scala 33:37]
  wire [2:0] _T_228 = _T_13 ? 3'h0 : _T_227; // @[Lookup.scala 33:37]
  wire [2:0] _T_229 = _T_11 ? 3'h0 : _T_228; // @[Lookup.scala 33:37]
  wire [2:0] _T_230 = _T_9 ? 3'h0 : _T_229; // @[Lookup.scala 33:37]
  wire [2:0] _T_231 = _T_7 ? 3'h0 : _T_230; // @[Lookup.scala 33:37]
  wire [2:0] _T_232 = _T_5 ? 3'h0 : _T_231; // @[Lookup.scala 33:37]
  wire [2:0] _T_233 = _T_3 ? 3'h0 : _T_232; // @[Lookup.scala 33:37]
  wire [5:0] _T_234 = _T_117 ? 6'h33 : 6'h0; // @[Lookup.scala 33:37]
  wire [5:0] _T_235 = _T_115 ? 6'h0 : _T_234; // @[Lookup.scala 33:37]
  wire [5:0] _T_236 = _T_113 ? 6'h32 : _T_235; // @[Lookup.scala 33:37]
  wire [5:0] _T_237 = _T_111 ? 6'h32 : _T_236; // @[Lookup.scala 33:37]
  wire [5:0] _T_238 = _T_109 ? 6'h31 : _T_237; // @[Lookup.scala 33:37]
  wire [5:0] _T_239 = _T_107 ? 6'h30 : _T_238; // @[Lookup.scala 33:37]
  wire [5:0] _T_240 = _T_105 ? 6'h2f : _T_239; // @[Lookup.scala 33:37]
  wire [5:0] _T_241 = _T_103 ? 6'h2e : _T_240; // @[Lookup.scala 33:37]
  wire [5:0] _T_242 = _T_101 ? 6'h2d : _T_241; // @[Lookup.scala 33:37]
  wire [5:0] _T_243 = _T_99 ? 6'h2c : _T_242; // @[Lookup.scala 33:37]
  wire [5:0] _T_244 = _T_97 ? 6'h2b : _T_243; // @[Lookup.scala 33:37]
  wire [5:0] _T_245 = _T_95 ? 6'h2a : _T_244; // @[Lookup.scala 33:37]
  wire [5:0] _T_246 = _T_93 ? 6'h29 : _T_245; // @[Lookup.scala 33:37]
  wire [5:0] _T_247 = _T_91 ? 6'h28 : _T_246; // @[Lookup.scala 33:37]
  wire [5:0] _T_248 = _T_89 ? 6'h26 : _T_247; // @[Lookup.scala 33:37]
  wire [5:0] _T_249 = _T_87 ? 6'h25 : _T_248; // @[Lookup.scala 33:37]
  wire [5:0] _T_250 = _T_85 ? 6'h24 : _T_249; // @[Lookup.scala 33:37]
  wire [5:0] _T_251 = _T_83 ? 6'h23 : _T_250; // @[Lookup.scala 33:37]
  wire [5:0] _T_252 = _T_81 ? 6'h22 : _T_251; // @[Lookup.scala 33:37]
  wire [5:0] _T_253 = _T_79 ? 6'h21 : _T_252; // @[Lookup.scala 33:37]
  wire [5:0] _T_254 = _T_77 ? 6'h20 : _T_253; // @[Lookup.scala 33:37]
  wire [5:0] _T_255 = _T_75 ? 6'h1f : _T_254; // @[Lookup.scala 33:37]
  wire [5:0] _T_256 = _T_73 ? 6'h1e : _T_255; // @[Lookup.scala 33:37]
  wire [5:0] _T_257 = _T_71 ? 6'h1d : _T_256; // @[Lookup.scala 33:37]
  wire [5:0] _T_258 = _T_69 ? 6'h1c : _T_257; // @[Lookup.scala 33:37]
  wire [5:0] _T_259 = _T_67 ? 6'h1b : _T_258; // @[Lookup.scala 33:37]
  wire [5:0] _T_260 = _T_65 ? 6'h1a : _T_259; // @[Lookup.scala 33:37]
  wire [5:0] _T_261 = _T_63 ? 6'h19 : _T_260; // @[Lookup.scala 33:37]
  wire [5:0] _T_262 = _T_61 ? 6'h18 : _T_261; // @[Lookup.scala 33:37]
  wire [5:0] _T_263 = _T_59 ? 6'h17 : _T_262; // @[Lookup.scala 33:37]
  wire [5:0] _T_264 = _T_57 ? 6'h10 : _T_263; // @[Lookup.scala 33:37]
  wire [5:0] _T_265 = _T_55 ? 6'h11 : _T_264; // @[Lookup.scala 33:37]
  wire [5:0] _T_266 = _T_53 ? 6'h16 : _T_265; // @[Lookup.scala 33:37]
  wire [5:0] _T_267 = _T_51 ? 6'h15 : _T_266; // @[Lookup.scala 33:37]
  wire [5:0] _T_268 = _T_49 ? 6'h11 : _T_267; // @[Lookup.scala 33:37]
  wire [5:0] _T_269 = _T_47 ? 6'h16 : _T_268; // @[Lookup.scala 33:37]
  wire [5:0] _T_270 = _T_45 ? 6'h15 : _T_269; // @[Lookup.scala 33:37]
  wire [5:0] _T_271 = _T_43 ? 6'h10 : _T_270; // @[Lookup.scala 33:37]
  wire [5:0] _T_272 = _T_41 ? 6'hf : _T_271; // @[Lookup.scala 33:37]
  wire [5:0] _T_273 = _T_39 ? 6'h0 : _T_272; // @[Lookup.scala 33:37]
  wire [5:0] _T_274 = _T_37 ? 6'hd : _T_273; // @[Lookup.scala 33:37]
  wire [5:0] _T_275 = _T_35 ? 6'h8 : _T_274; // @[Lookup.scala 33:37]
  wire [5:0] _T_276 = _T_33 ? 6'h7 : _T_275; // @[Lookup.scala 33:37]
  wire [5:0] _T_277 = _T_31 ? 6'h6 : _T_276; // @[Lookup.scala 33:37]
  wire [5:0] _T_278 = _T_29 ? 6'h5 : _T_277; // @[Lookup.scala 33:37]
  wire [5:0] _T_279 = _T_27 ? 6'h4 : _T_278; // @[Lookup.scala 33:37]
  wire [5:0] _T_280 = _T_25 ? 6'h3 : _T_279; // @[Lookup.scala 33:37]
  wire [5:0] _T_281 = _T_23 ? 6'h2 : _T_280; // @[Lookup.scala 33:37]
  wire [5:0] _T_282 = _T_21 ? 6'h1 : _T_281; // @[Lookup.scala 33:37]
  wire [5:0] _T_283 = _T_19 ? 6'h0 : _T_282; // @[Lookup.scala 33:37]
  wire [5:0] _T_284 = _T_17 ? 6'h6 : _T_283; // @[Lookup.scala 33:37]
  wire [5:0] _T_285 = _T_15 ? 6'h14 : _T_284; // @[Lookup.scala 33:37]
  wire [5:0] _T_286 = _T_13 ? 6'h7 : _T_285; // @[Lookup.scala 33:37]
  wire [5:0] _T_287 = _T_11 ? 6'h13 : _T_286; // @[Lookup.scala 33:37]
  wire [5:0] _T_288 = _T_9 ? 6'h4 : _T_287; // @[Lookup.scala 33:37]
  wire [5:0] _T_289 = _T_7 ? 6'h3 : _T_288; // @[Lookup.scala 33:37]
  wire [5:0] _T_290 = _T_5 ? 6'h2 : _T_289; // @[Lookup.scala 33:37]
  wire [5:0] _T_291 = _T_3 ? 6'h12 : _T_290; // @[Lookup.scala 33:37]
  wire  csri = io_op_type == 6'h2f | io_op_type == 6'h30 | io_op_type == 6'h31; // @[Decode.scala 30:63]
  wire  rs1_type = 3'h0 == instrType | (3'h7 == instrType | 3'h6 == instrType); // @[Mux.scala 80:57]
  wire  _io_rs2_type_T_1 = 3'h4 == instrType ? 1'h0 : 1'h1; // @[Mux.scala 80:57]
  wire  _io_rs2_type_T_5 = 3'h2 == instrType ? 1'h0 : 3'h5 == instrType | _io_rs2_type_T_1; // @[Mux.scala 80:57]
  wire  _io_rs2_type_T_7 = 3'h1 == instrType ? 1'h0 : _io_rs2_type_T_5; // @[Mux.scala 80:57]
  wire  _io_rs2_type_T_9 = 3'h6 == instrType ? 1'h0 : _io_rs2_type_T_7; // @[Mux.scala 80:57]
  wire  _io_rs2_type_T_11 = 3'h7 == instrType ? 1'h0 : _io_rs2_type_T_9; // @[Mux.scala 80:57]
  wire  _io_rs2_type_T_13 = 3'h0 == instrType ? 1'h0 : _io_rs2_type_T_11; // @[Mux.scala 80:57]
  wire [51:0] io_imm_hi = io_inst[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [11:0] io_imm_lo = io_inst[31:20]; // @[Decode.scala 58:45]
  wire [63:0] _io_imm_T_2 = {io_imm_hi,io_imm_lo}; // @[Cat.scala 30:58]
  wire [6:0] io_imm_hi_lo = io_inst[31:25]; // @[Decode.scala 59:45]
  wire [63:0] _io_imm_T_5 = {io_imm_hi,io_imm_hi_lo,io_inst[11:7]}; // @[Cat.scala 30:58]
  wire  io_imm_hi_hi_lo = io_inst[7]; // @[Decode.scala 60:45]
  wire [5:0] io_imm_hi_lo_1 = io_inst[30:25]; // @[Decode.scala 60:55]
  wire [3:0] io_imm_lo_hi = io_inst[11:8]; // @[Decode.scala 60:70]
  wire [63:0] _io_imm_T_8 = {io_imm_hi,io_imm_hi_hi_lo,io_imm_hi_lo_1,io_imm_lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire [31:0] io_imm_hi_hi_2 = io_inst[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [19:0] io_imm_hi_lo_2 = io_inst[31:12]; // @[Decode.scala 61:45]
  wire [63:0] _io_imm_T_11 = {io_imm_hi_hi_2,io_imm_hi_lo_2,12'h0}; // @[Cat.scala 30:58]
  wire [43:0] io_imm_hi_hi_hi_1 = io_inst[31] ? 44'hfffffffffff : 44'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_imm_hi_hi_lo_1 = io_inst[19:12]; // @[Decode.scala 62:45]
  wire  io_imm_hi_lo_3 = io_inst[20]; // @[Decode.scala 62:60]
  wire [9:0] io_imm_lo_hi_1 = io_inst[30:21]; // @[Decode.scala 62:71]
  wire [63:0] _io_imm_T_14 = {io_imm_hi_hi_hi_1,io_imm_hi_hi_lo_1,io_imm_hi_lo_3,io_imm_lo_hi_1,1'h0}; // @[Cat.scala 30:58]
  wire [63:0] _io_imm_T_16 = 3'h4 == instrType ? _io_imm_T_2 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_imm_T_18 = 3'h2 == instrType ? _io_imm_T_5 : _io_imm_T_16; // @[Mux.scala 80:57]
  wire [63:0] _io_imm_T_20 = 3'h1 == instrType ? _io_imm_T_8 : _io_imm_T_18; // @[Mux.scala 80:57]
  wire [63:0] _io_imm_T_22 = 3'h6 == instrType ? _io_imm_T_11 : _io_imm_T_20; // @[Mux.scala 80:57]
  wire [63:0] _io_csr_imm_T = {59'h0,io_inst[19:15]}; // @[Cat.scala 30:58]
  assign io_rs1_addr = instrType == 3'h6 | instrType == 3'h7 ? 5'h0 : io_inst[19:15]; // @[Decode.scala 27:21]
  assign io_rs1_type = csri ? 2'h2 : {{1'd0}, rs1_type}; // @[Decode.scala 46:21]
  assign io_rs2_addr = instrType == 3'h4 ? 5'h0 : io_inst[24:20]; // @[Decode.scala 28:21]
  assign io_rs2_type = {{1'd0}, _io_rs2_type_T_13}; // @[Mux.scala 80:57]
  assign io_rd_addr = instrType[2] ? io_inst[11:7] : 5'h0; // @[Decode.scala 34:20]
  assign io_rd_en = instrType[2]; // @[Decode.scala 31:50]
  assign io_op_type = _T_1 ? 6'h0 : _T_291; // @[Lookup.scala 33:37]
  assign io_fuType = _T_1 ? 3'h0 : _T_233; // @[Lookup.scala 33:37]
  assign io_imm = 3'h7 == instrType ? _io_imm_T_14 : _io_imm_T_22; // @[Mux.scala 80:57]
  assign io_csr_imm = csri ? _io_csr_imm_T : 64'h0; // @[Decode.scala 65:20]
endmodule
module ysyx_210340_RegFile(
  input         clock,
  input         reset,
  input  [31:0] io_pc,
  input  [4:0]  io_rs1_addr,
  input  [4:0]  io_rs2_addr,
  input  [1:0]  io_rs1_type,
  input  [1:0]  io_rs2_type,
  input  [4:0]  io_rd_addr,
  input         io_rd_en,
  input  [63:0] io_rd_data,
  input  [63:0] io_imm,
  input  [63:0] io_csr_imm,
  input         io_irq,
  output [63:0] io_rs1,
  output [63:0] io_rs2,
  output [63:0] io_src2
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] rf_0; // @[RegFile.scala 26:19]
  reg [63:0] rf_1; // @[RegFile.scala 26:19]
  reg [63:0] rf_2; // @[RegFile.scala 26:19]
  reg [63:0] rf_3; // @[RegFile.scala 26:19]
  reg [63:0] rf_4; // @[RegFile.scala 26:19]
  reg [63:0] rf_5; // @[RegFile.scala 26:19]
  reg [63:0] rf_6; // @[RegFile.scala 26:19]
  reg [63:0] rf_7; // @[RegFile.scala 26:19]
  reg [63:0] rf_8; // @[RegFile.scala 26:19]
  reg [63:0] rf_9; // @[RegFile.scala 26:19]
  reg [63:0] rf_10; // @[RegFile.scala 26:19]
  reg [63:0] rf_11; // @[RegFile.scala 26:19]
  reg [63:0] rf_12; // @[RegFile.scala 26:19]
  reg [63:0] rf_13; // @[RegFile.scala 26:19]
  reg [63:0] rf_14; // @[RegFile.scala 26:19]
  reg [63:0] rf_15; // @[RegFile.scala 26:19]
  reg [63:0] rf_16; // @[RegFile.scala 26:19]
  reg [63:0] rf_17; // @[RegFile.scala 26:19]
  reg [63:0] rf_18; // @[RegFile.scala 26:19]
  reg [63:0] rf_19; // @[RegFile.scala 26:19]
  reg [63:0] rf_20; // @[RegFile.scala 26:19]
  reg [63:0] rf_21; // @[RegFile.scala 26:19]
  reg [63:0] rf_22; // @[RegFile.scala 26:19]
  reg [63:0] rf_23; // @[RegFile.scala 26:19]
  reg [63:0] rf_24; // @[RegFile.scala 26:19]
  reg [63:0] rf_25; // @[RegFile.scala 26:19]
  reg [63:0] rf_26; // @[RegFile.scala 26:19]
  reg [63:0] rf_27; // @[RegFile.scala 26:19]
  reg [63:0] rf_28; // @[RegFile.scala 26:19]
  reg [63:0] rf_29; // @[RegFile.scala 26:19]
  reg [63:0] rf_30; // @[RegFile.scala 26:19]
  reg [63:0] rf_31; // @[RegFile.scala 26:19]
  wire [63:0] _GEN_1 = 5'h1 == io_rs1_addr ? rf_1 : rf_0; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_2 = 5'h2 == io_rs1_addr ? rf_2 : _GEN_1; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_3 = 5'h3 == io_rs1_addr ? rf_3 : _GEN_2; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_4 = 5'h4 == io_rs1_addr ? rf_4 : _GEN_3; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_5 = 5'h5 == io_rs1_addr ? rf_5 : _GEN_4; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_6 = 5'h6 == io_rs1_addr ? rf_6 : _GEN_5; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_7 = 5'h7 == io_rs1_addr ? rf_7 : _GEN_6; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_8 = 5'h8 == io_rs1_addr ? rf_8 : _GEN_7; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_9 = 5'h9 == io_rs1_addr ? rf_9 : _GEN_8; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_10 = 5'ha == io_rs1_addr ? rf_10 : _GEN_9; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_11 = 5'hb == io_rs1_addr ? rf_11 : _GEN_10; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_12 = 5'hc == io_rs1_addr ? rf_12 : _GEN_11; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_13 = 5'hd == io_rs1_addr ? rf_13 : _GEN_12; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_14 = 5'he == io_rs1_addr ? rf_14 : _GEN_13; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_15 = 5'hf == io_rs1_addr ? rf_15 : _GEN_14; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_16 = 5'h10 == io_rs1_addr ? rf_16 : _GEN_15; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_17 = 5'h11 == io_rs1_addr ? rf_17 : _GEN_16; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_18 = 5'h12 == io_rs1_addr ? rf_18 : _GEN_17; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_19 = 5'h13 == io_rs1_addr ? rf_19 : _GEN_18; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_20 = 5'h14 == io_rs1_addr ? rf_20 : _GEN_19; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_21 = 5'h15 == io_rs1_addr ? rf_21 : _GEN_20; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_22 = 5'h16 == io_rs1_addr ? rf_22 : _GEN_21; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_23 = 5'h17 == io_rs1_addr ? rf_23 : _GEN_22; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_24 = 5'h18 == io_rs1_addr ? rf_24 : _GEN_23; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_25 = 5'h19 == io_rs1_addr ? rf_25 : _GEN_24; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_26 = 5'h1a == io_rs1_addr ? rf_26 : _GEN_25; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_27 = 5'h1b == io_rs1_addr ? rf_27 : _GEN_26; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_28 = 5'h1c == io_rs1_addr ? rf_28 : _GEN_27; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_29 = 5'h1d == io_rs1_addr ? rf_29 : _GEN_28; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_30 = 5'h1e == io_rs1_addr ? rf_30 : _GEN_29; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_31 = 5'h1f == io_rs1_addr ? rf_31 : _GEN_30; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] rs1_data = io_rs1_addr == 5'h0 ? 64'h0 : _GEN_31; // @[RegFile.scala 27:36]
  wire [63:0] _GEN_33 = 5'h1 == io_rs2_addr ? rf_1 : rf_0; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_34 = 5'h2 == io_rs2_addr ? rf_2 : _GEN_33; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_35 = 5'h3 == io_rs2_addr ? rf_3 : _GEN_34; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_36 = 5'h4 == io_rs2_addr ? rf_4 : _GEN_35; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_37 = 5'h5 == io_rs2_addr ? rf_5 : _GEN_36; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_38 = 5'h6 == io_rs2_addr ? rf_6 : _GEN_37; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_39 = 5'h7 == io_rs2_addr ? rf_7 : _GEN_38; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_40 = 5'h8 == io_rs2_addr ? rf_8 : _GEN_39; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_41 = 5'h9 == io_rs2_addr ? rf_9 : _GEN_40; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_42 = 5'ha == io_rs2_addr ? rf_10 : _GEN_41; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_43 = 5'hb == io_rs2_addr ? rf_11 : _GEN_42; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_44 = 5'hc == io_rs2_addr ? rf_12 : _GEN_43; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_45 = 5'hd == io_rs2_addr ? rf_13 : _GEN_44; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_46 = 5'he == io_rs2_addr ? rf_14 : _GEN_45; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_47 = 5'hf == io_rs2_addr ? rf_15 : _GEN_46; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_48 = 5'h10 == io_rs2_addr ? rf_16 : _GEN_47; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_49 = 5'h11 == io_rs2_addr ? rf_17 : _GEN_48; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_50 = 5'h12 == io_rs2_addr ? rf_18 : _GEN_49; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_51 = 5'h13 == io_rs2_addr ? rf_19 : _GEN_50; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_52 = 5'h14 == io_rs2_addr ? rf_20 : _GEN_51; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_53 = 5'h15 == io_rs2_addr ? rf_21 : _GEN_52; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_54 = 5'h16 == io_rs2_addr ? rf_22 : _GEN_53; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_55 = 5'h17 == io_rs2_addr ? rf_23 : _GEN_54; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_56 = 5'h18 == io_rs2_addr ? rf_24 : _GEN_55; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_57 = 5'h19 == io_rs2_addr ? rf_25 : _GEN_56; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_58 = 5'h1a == io_rs2_addr ? rf_26 : _GEN_57; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_59 = 5'h1b == io_rs2_addr ? rf_27 : _GEN_58; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_60 = 5'h1c == io_rs2_addr ? rf_28 : _GEN_59; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_61 = 5'h1d == io_rs2_addr ? rf_29 : _GEN_60; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_62 = 5'h1e == io_rs2_addr ? rf_30 : _GEN_61; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] _GEN_63 = 5'h1f == io_rs2_addr ? rf_31 : _GEN_62; // @[RegFile.scala 27:36 RegFile.scala 27:36]
  wire [63:0] rs2_data = io_rs2_addr == 5'h0 ? 64'h0 : _GEN_63; // @[RegFile.scala 27:36]
  wire [63:0] _io_rs1_T_2 = io_rs1_type == 2'h2 ? io_csr_imm : rs1_data; // @[RegFile.scala 32:51]
  assign io_rs1 = io_rs1_type == 2'h1 ? {{32'd0}, io_pc} : _io_rs1_T_2; // @[RegFile.scala 32:16]
  assign io_rs2 = io_rs2_type == 2'h1 ? rs2_data : io_imm; // @[RegFile.scala 33:16]
  assign io_src2 = io_rs2_addr == 5'h0 ? 64'h0 : _GEN_63; // @[RegFile.scala 27:36]
  always @(posedge clock) begin
    if (reset) begin // @[RegFile.scala 26:19]
      rf_0 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h0 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_0 <= 64'h0;
        end else begin
          rf_0 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_1 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h1 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_1 <= 64'h0;
        end else begin
          rf_1 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_2 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h2 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_2 <= 64'h0;
        end else begin
          rf_2 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_3 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h3 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_3 <= 64'h0;
        end else begin
          rf_3 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_4 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h4 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_4 <= 64'h0;
        end else begin
          rf_4 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_5 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h5 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_5 <= 64'h0;
        end else begin
          rf_5 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_6 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h6 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_6 <= 64'h0;
        end else begin
          rf_6 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_7 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h7 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_7 <= 64'h0;
        end else begin
          rf_7 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_8 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h8 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_8 <= 64'h0;
        end else begin
          rf_8 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_9 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h9 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_9 <= 64'h0;
        end else begin
          rf_9 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_10 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'ha == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_10 <= 64'h0;
        end else begin
          rf_10 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_11 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'hb == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_11 <= 64'h0;
        end else begin
          rf_11 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_12 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'hc == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_12 <= 64'h0;
        end else begin
          rf_12 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_13 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'hd == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_13 <= 64'h0;
        end else begin
          rf_13 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_14 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'he == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_14 <= 64'h0;
        end else begin
          rf_14 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_15 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'hf == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_15 <= 64'h0;
        end else begin
          rf_15 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_16 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h10 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_16 <= 64'h0;
        end else begin
          rf_16 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_17 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h11 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_17 <= 64'h0;
        end else begin
          rf_17 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_18 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h12 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_18 <= 64'h0;
        end else begin
          rf_18 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_19 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h13 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_19 <= 64'h0;
        end else begin
          rf_19 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_20 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h14 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_20 <= 64'h0;
        end else begin
          rf_20 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_21 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h15 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_21 <= 64'h0;
        end else begin
          rf_21 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_22 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h16 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_22 <= 64'h0;
        end else begin
          rf_22 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_23 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h17 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_23 <= 64'h0;
        end else begin
          rf_23 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_24 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h18 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_24 <= 64'h0;
        end else begin
          rf_24 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_25 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h19 == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_25 <= 64'h0;
        end else begin
          rf_25 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_26 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h1a == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_26 <= 64'h0;
        end else begin
          rf_26 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_27 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h1b == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_27 <= 64'h0;
        end else begin
          rf_27 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_28 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h1c == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_28 <= 64'h0;
        end else begin
          rf_28 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_29 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h1d == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_29 <= 64'h0;
        end else begin
          rf_29 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_30 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h1e == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_30 <= 64'h0;
        end else begin
          rf_30 <= io_rd_data;
        end
      end
    end
    if (reset) begin // @[RegFile.scala 26:19]
      rf_31 <= 64'h0; // @[RegFile.scala 26:19]
    end else if (io_rd_en & ~io_irq) begin // @[RegFile.scala 36:30]
      if (5'h1f == io_rd_addr) begin // @[RegFile.scala 28:50]
        if (io_rd_addr == 5'h0) begin // @[RegFile.scala 28:56]
          rf_31 <= 64'h0;
        end else begin
          rf_31 <= io_rd_data;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  rf_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  rf_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  rf_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  rf_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  rf_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  rf_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  rf_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  rf_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  rf_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  rf_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  rf_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  rf_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  rf_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  rf_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  rf_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  rf_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  rf_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  rf_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  rf_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  rf_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  rf_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  rf_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  rf_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  rf_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  rf_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  rf_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  rf_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  rf_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  rf_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  rf_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  rf_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  rf_31 = _RAND_31[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210340_Execution(
  input  [31:0] io_pc,
  input  [5:0]  io_op_type,
  input  [63:0] io_rs1,
  input  [63:0] io_rs2,
  input  [63:0] io_src2,
  input  [2:0]  io_fuType,
  input  [63:0] io_imm,
  input  [31:0] io_csr_Jmp_addr,
  input         io_csr_Jmp_en,
  input  [63:0] io_csr_data,
  output        io_br_en,
  output [31:0] io_br_addr,
  output [63:0] io_rd_data,
  output        fence_i_0
);
  wire  fence_i = io_fuType == 3'h4; // @[Execution.scala 25:28]
  wire [4:0] aluOut_shamt = io_rs2[4:0]; // @[Execution.scala 29:20]
  wire [5:0] aluOut_shamt64 = io_imm[5:0]; // @[Execution.scala 30:22]
  wire [31:0] _aluOut_sraw_T_1 = io_rs1[31:0]; // @[Execution.scala 31:29]
  wire [31:0] aluOut_sraw = $signed(_aluOut_sraw_T_1) >>> aluOut_shamt; // @[Execution.scala 31:46]
  wire [63:0] _aluOut_T_1 = io_rs1 + io_rs2; // @[Execution.scala 33:24]
  wire [126:0] _GEN_4 = {{63'd0}, io_rs1}; // @[Execution.scala 34:23]
  wire [126:0] _aluOut_T_3 = _GEN_4 << io_rs2[5:0]; // @[Execution.scala 34:23]
  wire [126:0] _aluOut_T_4 = _GEN_4 << aluOut_shamt64; // @[Execution.scala 35:23]
  wire  _aluOut_T_7 = $signed(io_rs1) < $signed(io_rs2); // @[Execution.scala 36:31]
  wire  _aluOut_T_8 = io_rs1 < io_rs2; // @[Execution.scala 37:24]
  wire [63:0] _aluOut_T_9 = io_rs1 ^ io_rs2; // @[Execution.scala 38:24]
  wire [63:0] _aluOut_T_10 = io_rs1 >> aluOut_shamt; // @[Execution.scala 39:24]
  wire [63:0] _aluOut_T_11 = io_rs1 >> aluOut_shamt64; // @[Execution.scala 40:24]
  wire [63:0] _aluOut_T_12 = io_rs1 | io_rs2; // @[Execution.scala 41:24]
  wire [63:0] _aluOut_T_13 = io_rs1 & io_rs2; // @[Execution.scala 42:24]
  wire [63:0] _aluOut_T_15 = io_rs1 - io_rs2; // @[Execution.scala 43:24]
  wire [63:0] _aluOut_T_18 = $signed(io_rs1) >>> aluOut_shamt; // @[Execution.scala 45:41]
  wire [63:0] _aluOut_T_21 = $signed(io_rs1) >>> aluOut_shamt64; // @[Execution.scala 46:43]
  wire [31:0] aluOut_hi = _aluOut_T_1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] aluOut_lo = _aluOut_T_1[31:0]; // @[Execution.scala 47:60]
  wire [63:0] _aluOut_T_28 = {aluOut_hi,aluOut_lo}; // @[Cat.scala 30:58]
  wire [31:0] aluOut_hi_1 = aluOut_sraw[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _aluOut_T_31 = {aluOut_hi_1,aluOut_sraw}; // @[Cat.scala 30:58]
  wire [62:0] _GEN_6 = {{31'd0}, io_rs1[31:0]}; // @[Execution.scala 49:44]
  wire [62:0] _aluOut_T_33 = _GEN_6 << aluOut_shamt; // @[Execution.scala 49:44]
  wire [31:0] aluOut_hi_2 = _aluOut_T_33[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] aluOut_lo_2 = _aluOut_T_33[31:0]; // @[Execution.scala 49:80]
  wire [63:0] _aluOut_T_38 = {aluOut_hi_2,aluOut_lo_2}; // @[Cat.scala 30:58]
  wire [31:0] _aluOut_T_40 = io_rs1[31:0] >> aluOut_shamt; // @[Execution.scala 50:44]
  wire [31:0] aluOut_hi_3 = _aluOut_T_40[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _aluOut_T_45 = {aluOut_hi_3,_aluOut_T_40}; // @[Cat.scala 30:58]
  wire [31:0] aluOut_hi_4 = _aluOut_T_15[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] aluOut_lo_4 = _aluOut_T_15[31:0]; // @[Execution.scala 51:60]
  wire [63:0] _aluOut_T_52 = {aluOut_hi_4,aluOut_lo_4}; // @[Cat.scala 30:58]
  wire [63:0] _aluOut_T_54 = 6'h0 == io_op_type ? _aluOut_T_1 : 64'h0; // @[Mux.scala 80:57]
  wire [126:0] _aluOut_T_56 = 6'h1 == io_op_type ? _aluOut_T_3 : {{63'd0}, _aluOut_T_54}; // @[Mux.scala 80:57]
  wire [126:0] _aluOut_T_58 = 6'h12 == io_op_type ? _aluOut_T_4 : _aluOut_T_56; // @[Mux.scala 80:57]
  wire [126:0] _aluOut_T_60 = 6'h2 == io_op_type ? {{126'd0}, _aluOut_T_7} : _aluOut_T_58; // @[Mux.scala 80:57]
  wire [126:0] _aluOut_T_62 = 6'h3 == io_op_type ? {{126'd0}, _aluOut_T_8} : _aluOut_T_60; // @[Mux.scala 80:57]
  wire [126:0] _aluOut_T_64 = 6'h4 == io_op_type ? {{63'd0}, _aluOut_T_9} : _aluOut_T_62; // @[Mux.scala 80:57]
  wire [126:0] _aluOut_T_66 = 6'h5 == io_op_type ? {{63'd0}, _aluOut_T_10} : _aluOut_T_64; // @[Mux.scala 80:57]
  wire [126:0] _aluOut_T_68 = 6'h13 == io_op_type ? {{63'd0}, _aluOut_T_11} : _aluOut_T_66; // @[Mux.scala 80:57]
  wire [126:0] _aluOut_T_70 = 6'h6 == io_op_type ? {{63'd0}, _aluOut_T_12} : _aluOut_T_68; // @[Mux.scala 80:57]
  wire [126:0] _aluOut_T_72 = 6'h7 == io_op_type ? {{63'd0}, _aluOut_T_13} : _aluOut_T_70; // @[Mux.scala 80:57]
  wire [126:0] _aluOut_T_74 = 6'h8 == io_op_type ? {{63'd0}, _aluOut_T_15} : _aluOut_T_72; // @[Mux.scala 80:57]
  wire [126:0] _aluOut_T_76 = 6'hf == io_op_type ? {{63'd0}, io_rs2} : _aluOut_T_74; // @[Mux.scala 80:57]
  wire [126:0] _aluOut_T_78 = 6'hd == io_op_type ? {{63'd0}, _aluOut_T_18} : _aluOut_T_76; // @[Mux.scala 80:57]
  wire [126:0] _aluOut_T_80 = 6'h14 == io_op_type ? {{63'd0}, _aluOut_T_21} : _aluOut_T_78; // @[Mux.scala 80:57]
  wire [126:0] _aluOut_T_82 = 6'h10 == io_op_type ? {{63'd0}, _aluOut_T_28} : _aluOut_T_80; // @[Mux.scala 80:57]
  wire [126:0] _aluOut_T_84 = 6'h11 == io_op_type ? {{63'd0}, _aluOut_T_31} : _aluOut_T_82; // @[Mux.scala 80:57]
  wire [126:0] _aluOut_T_86 = 6'h15 == io_op_type ? {{63'd0}, _aluOut_T_38} : _aluOut_T_84; // @[Mux.scala 80:57]
  wire [126:0] _aluOut_T_88 = 6'h16 == io_op_type ? {{63'd0}, _aluOut_T_45} : _aluOut_T_86; // @[Mux.scala 80:57]
  wire [126:0] aluOut = 6'h17 == io_op_type ? {{63'd0}, _aluOut_T_52} : _aluOut_T_88; // @[Mux.scala 80:57]
  wire  _jmp_en_T = io_fuType == 3'h1; // @[Execution.scala 69:35]
  wire  _jmp_en_T_1 = io_rs1 == io_src2; // @[Execution.scala 57:23]
  wire  _jmp_en_T_2 = io_rs1 != io_src2; // @[Execution.scala 58:23]
  wire  _jmp_en_T_5 = $signed(io_rs1) < $signed(io_src2); // @[Execution.scala 59:31]
  wire  _jmp_en_T_8 = $signed(io_rs1) >= $signed(io_src2); // @[Execution.scala 60:30]
  wire  _jmp_en_T_9 = io_rs1 < io_src2; // @[Execution.scala 61:24]
  wire  _jmp_en_T_10 = io_rs1 >= io_src2; // @[Execution.scala 62:24]
  wire  _jmp_en_T_14 = 6'h1b == io_op_type ? _jmp_en_T_2 : 6'h1a == io_op_type & _jmp_en_T_1; // @[Mux.scala 80:57]
  wire  _jmp_en_T_16 = 6'h1c == io_op_type ? _jmp_en_T_5 : _jmp_en_T_14; // @[Mux.scala 80:57]
  wire  _jmp_en_T_18 = 6'h1d == io_op_type ? _jmp_en_T_8 : _jmp_en_T_16; // @[Mux.scala 80:57]
  wire  _jmp_en_T_20 = 6'h1e == io_op_type ? _jmp_en_T_9 : _jmp_en_T_18; // @[Mux.scala 80:57]
  wire  _jmp_en_T_22 = 6'h1f == io_op_type ? _jmp_en_T_10 : _jmp_en_T_20; // @[Mux.scala 80:57]
  wire  _jmp_en_T_26 = 6'h19 == io_op_type | (6'h18 == io_op_type | _jmp_en_T_22); // @[Mux.scala 80:57]
  wire  jmp_en = _jmp_en_T & _jmp_en_T_26; // @[Execution.scala 56:11]
  wire [63:0] _GEN_8 = {{32'd0}, io_pc}; // @[Execution.scala 70:69]
  wire [63:0] _jmp_addr_T_4 = _GEN_8 + io_rs2; // @[Execution.scala 70:69]
  wire [63:0] jmp_addr = io_op_type == 6'h19 ? _aluOut_T_1 : _jmp_addr_T_4; // @[Execution.scala 70:21]
  wire [31:0] _io_rd_data_T_1 = io_pc + 32'h4; // @[Execution.scala 74:21]
  wire [126:0] _io_rd_data_T_3 = 3'h0 == io_fuType ? aluOut : 127'h0; // @[Mux.scala 80:57]
  wire [126:0] _io_rd_data_T_5 = 3'h1 == io_fuType ? {{95'd0}, _io_rd_data_T_1} : _io_rd_data_T_3; // @[Mux.scala 80:57]
  wire [126:0] _io_rd_data_T_7 = 3'h3 == io_fuType ? {{63'd0}, io_csr_data} : _io_rd_data_T_5; // @[Mux.scala 80:57]
  wire [126:0] _io_rd_data_T_9 = 3'h4 == io_fuType ? 127'h0 : _io_rd_data_T_7; // @[Mux.scala 80:57]
  wire  _GEN_0 = io_csr_Jmp_en ? io_csr_Jmp_en : jmp_en; // @[Execution.scala 83:29 Execution.scala 84:14 Execution.scala 87:14]
  wire [63:0] _GEN_1 = io_csr_Jmp_en ? {{32'd0}, io_csr_Jmp_addr} : jmp_addr; // @[Execution.scala 83:29 Execution.scala 85:16 Execution.scala 88:16]
  wire [63:0] _GEN_3 = fence_i ? {{32'd0}, _io_rd_data_T_1} : _GEN_1; // @[Execution.scala 79:19 Execution.scala 81:16]
  assign io_br_en = fence_i | _GEN_0; // @[Execution.scala 79:19 Execution.scala 80:14]
  assign io_br_addr = _GEN_3[31:0];
  assign io_rd_data = _io_rd_data_T_9[63:0]; // @[Execution.scala 72:13]
  assign fence_i_0 = fence_i;
endmodule
module ysyx_210340_PipelineReg_1(
  input         clock,
  input         reset,
  input  [31:0] io_in_pc,
  input         io_in_br_en,
  input  [31:0] io_in_br_addr,
  input  [5:0]  io_in_op_type,
  input  [2:0]  io_in_fuType,
  input  [63:0] io_in_rs1,
  input  [63:0] io_in_rs2,
  input  [4:0]  io_in_rd_addr,
  input  [63:0] io_in_src2,
  input         io_in_rd_en,
  input         io_in_imem_hs,
  input  [63:0] io_in_rd_data,
  output [31:0] io_out_pc,
  output        io_out_br_en,
  output [31:0] io_out_br_addr,
  output [5:0]  io_out_op_type,
  output [2:0]  io_out_fuType,
  output [63:0] io_out_rs1,
  output [63:0] io_out_rs2,
  output [4:0]  io_out_rd_addr,
  output [63:0] io_out_src2,
  output        io_out_rd_en,
  output        io_out_imem_hs,
  output [63:0] io_out_rd_data,
  input         io_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_pc; // @[PipelineReg.scala 60:20]
  reg  reg_br_en; // @[PipelineReg.scala 60:20]
  reg [31:0] reg_br_addr; // @[PipelineReg.scala 60:20]
  reg [5:0] reg_op_type; // @[PipelineReg.scala 60:20]
  reg [2:0] reg_fuType; // @[PipelineReg.scala 60:20]
  reg [63:0] reg_rs1; // @[PipelineReg.scala 60:20]
  reg [63:0] reg_rs2; // @[PipelineReg.scala 60:20]
  reg [4:0] reg_rd_addr; // @[PipelineReg.scala 60:20]
  reg [63:0] reg_src2; // @[PipelineReg.scala 60:20]
  reg  reg_rd_en; // @[PipelineReg.scala 60:20]
  reg  reg_imem_hs; // @[PipelineReg.scala 60:20]
  reg [63:0] reg_rd_data; // @[PipelineReg.scala 60:20]
  assign io_out_pc = reg_pc; // @[PipelineReg.scala 68:10]
  assign io_out_br_en = reg_br_en; // @[PipelineReg.scala 68:10]
  assign io_out_br_addr = reg_br_addr; // @[PipelineReg.scala 68:10]
  assign io_out_op_type = reg_op_type; // @[PipelineReg.scala 68:10]
  assign io_out_fuType = reg_fuType; // @[PipelineReg.scala 68:10]
  assign io_out_rs1 = reg_rs1; // @[PipelineReg.scala 68:10]
  assign io_out_rs2 = reg_rs2; // @[PipelineReg.scala 68:10]
  assign io_out_rd_addr = reg_rd_addr; // @[PipelineReg.scala 68:10]
  assign io_out_src2 = reg_src2; // @[PipelineReg.scala 68:10]
  assign io_out_rd_en = reg_rd_en; // @[PipelineReg.scala 68:10]
  assign io_out_imem_hs = reg_imem_hs; // @[PipelineReg.scala 68:10]
  assign io_out_rd_data = reg_rd_data; // @[PipelineReg.scala 68:10]
  always @(posedge clock) begin
    if (reset) begin // @[PipelineReg.scala 60:20]
      reg_pc <= 32'h0; // @[PipelineReg.scala 60:20]
    end else if (~io_stall) begin // @[PipelineReg.scala 64:27]
      reg_pc <= io_in_pc; // @[PipelineReg.scala 65:9]
    end
    if (reset) begin // @[PipelineReg.scala 60:20]
      reg_br_en <= 1'h0; // @[PipelineReg.scala 60:20]
    end else if (~io_stall) begin // @[PipelineReg.scala 64:27]
      reg_br_en <= io_in_br_en; // @[PipelineReg.scala 65:9]
    end
    if (reset) begin // @[PipelineReg.scala 60:20]
      reg_br_addr <= 32'h0; // @[PipelineReg.scala 60:20]
    end else if (~io_stall) begin // @[PipelineReg.scala 64:27]
      reg_br_addr <= io_in_br_addr; // @[PipelineReg.scala 65:9]
    end
    if (reset) begin // @[PipelineReg.scala 60:20]
      reg_op_type <= 6'h0; // @[PipelineReg.scala 60:20]
    end else if (~io_stall) begin // @[PipelineReg.scala 64:27]
      reg_op_type <= io_in_op_type; // @[PipelineReg.scala 65:9]
    end
    if (reset) begin // @[PipelineReg.scala 60:20]
      reg_fuType <= 3'h0; // @[PipelineReg.scala 60:20]
    end else if (~io_stall) begin // @[PipelineReg.scala 64:27]
      reg_fuType <= io_in_fuType; // @[PipelineReg.scala 65:9]
    end
    if (reset) begin // @[PipelineReg.scala 60:20]
      reg_rs1 <= 64'h0; // @[PipelineReg.scala 60:20]
    end else if (~io_stall) begin // @[PipelineReg.scala 64:27]
      reg_rs1 <= io_in_rs1; // @[PipelineReg.scala 65:9]
    end
    if (reset) begin // @[PipelineReg.scala 60:20]
      reg_rs2 <= 64'h0; // @[PipelineReg.scala 60:20]
    end else if (~io_stall) begin // @[PipelineReg.scala 64:27]
      reg_rs2 <= io_in_rs2; // @[PipelineReg.scala 65:9]
    end
    if (reset) begin // @[PipelineReg.scala 60:20]
      reg_rd_addr <= 5'h0; // @[PipelineReg.scala 60:20]
    end else if (~io_stall) begin // @[PipelineReg.scala 64:27]
      reg_rd_addr <= io_in_rd_addr; // @[PipelineReg.scala 65:9]
    end
    if (reset) begin // @[PipelineReg.scala 60:20]
      reg_src2 <= 64'h0; // @[PipelineReg.scala 60:20]
    end else if (~io_stall) begin // @[PipelineReg.scala 64:27]
      reg_src2 <= io_in_src2; // @[PipelineReg.scala 65:9]
    end
    if (reset) begin // @[PipelineReg.scala 60:20]
      reg_rd_en <= 1'h0; // @[PipelineReg.scala 60:20]
    end else if (~io_stall) begin // @[PipelineReg.scala 64:27]
      reg_rd_en <= io_in_rd_en; // @[PipelineReg.scala 65:9]
    end
    if (reset) begin // @[PipelineReg.scala 60:20]
      reg_imem_hs <= 1'h0; // @[PipelineReg.scala 60:20]
    end else if (~io_stall) begin // @[PipelineReg.scala 64:27]
      reg_imem_hs <= io_in_imem_hs; // @[PipelineReg.scala 65:9]
    end
    if (reset) begin // @[PipelineReg.scala 60:20]
      reg_rd_data <= 64'h0; // @[PipelineReg.scala 60:20]
    end else if (~io_stall) begin // @[PipelineReg.scala 64:27]
      reg_rd_data <= io_in_rd_data; // @[PipelineReg.scala 65:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_br_en = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  reg_br_addr = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_op_type = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  reg_fuType = _RAND_4[2:0];
  _RAND_5 = {2{`RANDOM}};
  reg_rs1 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  reg_rs2 = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  reg_rd_addr = _RAND_7[4:0];
  _RAND_8 = {2{`RANDOM}};
  reg_src2 = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  reg_rd_en = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  reg_imem_hs = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  reg_rd_data = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210340_Mem(
  input         clock,
  input         reset,
  input  [31:0] io_pc,
  input  [5:0]  io_op_type,
  input  [63:0] io_rs1,
  input  [63:0] io_rs2,
  input  [63:0] io_src2,
  input  [2:0]  io_fuType,
  input         io_irq,
  output        io_mem_en,
  output [63:0] io_rd_data,
  output        io_busy,
  output        io_dmem_hs,
  output        io_resp_success,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [31:0] io_dmem_req_bits_addr,
  output        io_dmem_req_bits_ren,
  output [63:0] io_dmem_req_bits_wdata,
  output [7:0]  io_dmem_req_bits_wmask,
  output        io_dmem_req_bits_wen,
  output [1:0]  io_dmem_req_bits_size,
  output        io_dmem_resp_ready,
  input         io_dmem_resp_valid,
  input  [63:0] io_dmem_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[Mem.scala 26:22]
  wire [63:0] _addr_T_1 = io_rs1 + io_rs2; // @[Mem.scala 31:22]
  wire [31:0] addr = _addr_T_1[31:0]; // @[Mem.scala 31:31]
  reg [31:0] reg_addr; // @[Mem.scala 34:25]
  wire [2:0] reg_addr_offset = reg_addr[2:0]; // @[Mem.scala 35:33]
  reg [63:0] reg_wdata; // @[Mem.scala 36:26]
  wire  mem_en = io_fuType == 3'h2; // @[Mem.scala 38:27]
  wire  mem_ren = mem_en & ~io_op_type[3]; // @[Mem.scala 39:37]
  wire  mem_wen = mem_en & io_op_type[3]; // @[Mem.scala 40:37]
  wire  mmio = ~addr[31] & io_pc != 32'h0; // @[Mem.scala 43:33]
  wire [7:0] _mask_T_1 = 3'h1 == reg_addr_offset ? 8'hfe : 8'hff; // @[Mux.scala 80:57]
  wire [7:0] _mask_T_3 = 3'h2 == reg_addr_offset ? 8'hfc : _mask_T_1; // @[Mux.scala 80:57]
  wire [7:0] _mask_T_5 = 3'h3 == reg_addr_offset ? 8'hf8 : _mask_T_3; // @[Mux.scala 80:57]
  wire [7:0] _mask_T_7 = 3'h4 == reg_addr_offset ? 8'hf0 : _mask_T_5; // @[Mux.scala 80:57]
  wire [7:0] _mask_T_9 = 3'h5 == reg_addr_offset ? 8'he0 : _mask_T_7; // @[Mux.scala 80:57]
  wire [7:0] _mask_T_11 = 3'h6 == reg_addr_offset ? 8'hc0 : _mask_T_9; // @[Mux.scala 80:57]
  wire [7:0] mask = 3'h7 == reg_addr_offset ? 8'h80 : _mask_T_11; // @[Mux.scala 80:57]
  wire [1:0] _wmask_T_3 = 6'h29 == io_op_type ? 2'h3 : {{1'd0}, 6'h28 == io_op_type}; // @[Mux.scala 80:57]
  wire [3:0] _wmask_T_5 = 6'h2a == io_op_type ? 4'hf : {{2'd0}, _wmask_T_3}; // @[Mux.scala 80:57]
  wire [7:0] wmask = 6'h2b == io_op_type ? 8'hff : {{4'd0}, _wmask_T_5}; // @[Mux.scala 80:57]
  wire [1:0] _inst_size_T_5 = 6'h2a == io_op_type ? 2'h2 : {{1'd0}, 6'h29 == io_op_type}; // @[Mux.scala 80:57]
  wire [1:0] _inst_size_T_7 = 6'h2b == io_op_type ? 2'h3 : _inst_size_T_5; // @[Mux.scala 80:57]
  wire [1:0] _inst_size_T_9 = 6'h20 == io_op_type ? 2'h0 : _inst_size_T_7; // @[Mux.scala 80:57]
  wire [1:0] _inst_size_T_11 = 6'h21 == io_op_type ? 2'h1 : _inst_size_T_9; // @[Mux.scala 80:57]
  wire [1:0] _inst_size_T_13 = 6'h22 == io_op_type ? 2'h2 : _inst_size_T_11; // @[Mux.scala 80:57]
  wire [1:0] _inst_size_T_15 = 6'h23 == io_op_type ? 2'h3 : _inst_size_T_13; // @[Mux.scala 80:57]
  wire [1:0] _inst_size_T_17 = 6'h24 == io_op_type ? 2'h0 : _inst_size_T_15; // @[Mux.scala 80:57]
  wire [1:0] _inst_size_T_19 = 6'h25 == io_op_type ? 2'h1 : _inst_size_T_17; // @[Mux.scala 80:57]
  wire [1:0] inst_size = 6'h26 == io_op_type ? 2'h2 : _inst_size_T_19; // @[Mux.scala 80:57]
  wire [28:0] io_dmem_req_bits_addr_hi = reg_addr[31:3]; // @[Mem.scala 78:48]
  wire [31:0] _io_dmem_req_bits_addr_T = {io_dmem_req_bits_addr_hi,3'h0}; // @[Cat.scala 30:58]
  wire [5:0] _io_dmem_req_bits_wdata_T = {reg_addr_offset, 3'h0}; // @[Mem.scala 80:52]
  wire [126:0] _GEN_22 = {{63'd0}, reg_wdata}; // @[Mem.scala 80:32]
  wire [126:0] _io_dmem_req_bits_wdata_T_1 = _GEN_22 << _io_dmem_req_bits_wdata_T; // @[Mem.scala 80:32]
  wire [14:0] _GEN_23 = {{7'd0}, wmask}; // @[Mem.scala 81:36]
  wire [14:0] _io_dmem_req_bits_wmask_T = _GEN_23 << reg_addr_offset; // @[Mem.scala 81:36]
  wire  _io_dmem_req_valid_T = state == 3'h1; // @[Mem.scala 85:23]
  wire  _io_dmem_req_valid_T_3 = ~io_irq; // @[Mem.scala 85:61]
  wire  _io_dmem_resp_ready_T = state == 3'h2; // @[Mem.scala 87:24]
  wire  _io_dmem_resp_ready_T_1 = state == 3'h3; // @[Mem.scala 87:48]
  reg [63:0] ram_rdata; // @[Mem.scala 89:26]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = io_dmem_req_ready & io_dmem_req_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_3 = mem_wen & _T_4 ? 3'h3 : state; // @[Mem.scala 110:43 Mem.scala 111:15 Mem.scala 26:22]
  wire [2:0] _GEN_4 = mem_ren & _T_4 ? 3'h2 : _GEN_3; // @[Mem.scala 108:43 Mem.scala 109:15]
  wire  _T_8 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [63:0] _ram_rdata_T_1 = io_dmem_resp_bits_rdata >> _io_dmem_req_bits_wdata_T; // @[Mem.scala 116:38]
  wire [63:0] _GEN_6 = io_resp_success ? _ram_rdata_T_1 : ram_rdata; // @[Mem.scala 115:30 Mem.scala 116:19 Mem.scala 89:26]
  wire [2:0] _GEN_7 = io_resp_success ? 3'h4 : state; // @[Mem.scala 115:30 Mem.scala 118:15 Mem.scala 26:22]
  wire  _T_9 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_10 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_8 = _T_10 ? 3'h0 : state; // @[Conditional.scala 39:67 Mem.scala 127:13 Mem.scala 26:22]
  wire [31:0] _GEN_9 = _T_10 ? 32'h0 : reg_addr; // @[Conditional.scala 39:67 Mem.scala 128:16 Mem.scala 34:25]
  wire [2:0] _GEN_10 = _T_9 ? _GEN_7 : _GEN_8; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_11 = _T_9 ? reg_addr : _GEN_9; // @[Conditional.scala 39:67 Mem.scala 34:25]
  wire [55:0] load_out_hi = ram_rdata[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [7:0] load_out_lo = ram_rdata[7:0]; // @[Mem.scala 135:55]
  wire [63:0] _load_out_T_2 = {load_out_hi,load_out_lo}; // @[Cat.scala 30:58]
  wire [47:0] load_out_hi_1 = ram_rdata[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [15:0] load_out_lo_1 = ram_rdata[15:0]; // @[Mem.scala 136:56]
  wire [63:0] _load_out_T_5 = {load_out_hi_1,load_out_lo_1}; // @[Cat.scala 30:58]
  wire [31:0] load_out_hi_2 = ram_rdata[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] load_out_lo_2 = ram_rdata[31:0]; // @[Mem.scala 137:56]
  wire [63:0] _load_out_T_8 = {load_out_hi_2,load_out_lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _load_out_T_9 = {56'h0,load_out_lo}; // @[Cat.scala 30:58]
  wire [63:0] _load_out_T_10 = {48'h0,load_out_lo_1}; // @[Cat.scala 30:58]
  wire [63:0] _load_out_T_11 = {32'h0,load_out_lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _load_out_T_13 = 6'h20 == io_op_type ? _load_out_T_2 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _load_out_T_15 = 6'h21 == io_op_type ? _load_out_T_5 : _load_out_T_13; // @[Mux.scala 80:57]
  wire [63:0] _load_out_T_17 = 6'h22 == io_op_type ? _load_out_T_8 : _load_out_T_15; // @[Mux.scala 80:57]
  wire [63:0] _load_out_T_19 = 6'h23 == io_op_type ? ram_rdata : _load_out_T_17; // @[Mux.scala 80:57]
  wire [63:0] _load_out_T_21 = 6'h24 == io_op_type ? _load_out_T_9 : _load_out_T_19; // @[Mux.scala 80:57]
  wire [63:0] _load_out_T_23 = 6'h25 == io_op_type ? _load_out_T_10 : _load_out_T_21; // @[Mux.scala 80:57]
  wire [63:0] load_out = 6'h26 == io_op_type ? _load_out_T_11 : _load_out_T_23; // @[Mux.scala 80:57]
  wire  _io_busy_T_5 = state == 3'h0 & mem_en | _io_dmem_req_valid_T | _io_dmem_resp_ready_T; // @[Mem.scala 158:66]
  assign io_mem_en = io_fuType == 3'h2; // @[Mem.scala 38:27]
  assign io_rd_data = state == 3'h4 ? load_out : 64'h0; // @[Mem.scala 157:20]
  assign io_busy = _io_busy_T_5 | _io_dmem_resp_ready_T_1; // @[Mem.scala 159:35]
  assign io_dmem_hs = io_dmem_resp_ready & io_dmem_resp_valid; // @[Mem.scala 95:28]
  assign io_resp_success = io_dmem_resp_ready & io_dmem_resp_valid; // @[Decoupled.scala 40:37]
  assign io_dmem_req_valid = state == 3'h1 & (mem_ren | mem_wen) & ~io_irq; // @[Mem.scala 85:58]
  assign io_dmem_req_bits_addr = mmio ? addr : _io_dmem_req_bits_addr_T; // @[Mem.scala 78:23]
  assign io_dmem_req_bits_ren = mem_en & ~io_op_type[3]; // @[Mem.scala 39:37]
  assign io_dmem_req_bits_wdata = _io_dmem_req_bits_wdata_T_1[63:0]; // @[Mem.scala 80:58]
  assign io_dmem_req_bits_wmask = mask & _io_dmem_req_bits_wmask_T[7:0]; // @[Mem.scala 81:26]
  assign io_dmem_req_bits_wen = mem_en & io_op_type[3]; // @[Mem.scala 40:37]
  assign io_dmem_req_bits_size = mmio ? inst_size : 2'h3; // @[Mem.scala 83:23]
  assign io_dmem_resp_ready = state == 3'h2 | state == 3'h3; // @[Mem.scala 87:38]
  always @(posedge clock) begin
    if (reset) begin // @[Mem.scala 26:22]
      state <= 3'h0; // @[Mem.scala 26:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (mem_en & _io_dmem_req_valid_T_3) begin // @[Mem.scala 99:31]
        state <= 3'h1; // @[Mem.scala 100:15]
      end
    end else if (_T_3) begin // @[Conditional.scala 39:67]
      if (io_irq) begin // @[Mem.scala 106:21]
        state <= 3'h0; // @[Mem.scala 107:15]
      end else begin
        state <= _GEN_4;
      end
    end else if (_T_8) begin // @[Conditional.scala 39:67]
      state <= _GEN_7;
    end else begin
      state <= _GEN_10;
    end
    if (reset) begin // @[Mem.scala 34:25]
      reg_addr <= 32'h0; // @[Mem.scala 34:25]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (mem_en & _io_dmem_req_valid_T_3) begin // @[Mem.scala 99:31]
        reg_addr <= addr; // @[Mem.scala 101:18]
      end
    end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
      if (!(_T_8)) begin // @[Conditional.scala 39:67]
        reg_addr <= _GEN_11;
      end
    end
    if (reset) begin // @[Mem.scala 36:26]
      reg_wdata <= 64'h0; // @[Mem.scala 36:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (mem_en & _io_dmem_req_valid_T_3) begin // @[Mem.scala 99:31]
        reg_wdata <= io_src2; // @[Mem.scala 102:19]
      end
    end
    if (reset) begin // @[Mem.scala 89:26]
      ram_rdata <= 64'h0; // @[Mem.scala 89:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_3)) begin // @[Conditional.scala 39:67]
        if (_T_8) begin // @[Conditional.scala 39:67]
          ram_rdata <= _GEN_6;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  reg_addr = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  reg_wdata = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  ram_rdata = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210340_CSR(
  input         clock,
  input         reset,
  input  [31:0] io_pc,
  input  [2:0]  io_fuType,
  input  [5:0]  io_op_type,
  input  [63:0] io_rs1,
  input  [63:0] io_rs2,
  input         io_if_valid,
  input         io_mem_en,
  input         io_mem_valid,
  output [31:0] io_csr_Jmp_addr,
  output        io_csr_Jmp_en,
  output [63:0] io_csr_data,
  output        io_irq,
  input         mtip_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtvec; // @[CSR.scala 25:26]
  reg [63:0] mcause; // @[CSR.scala 26:26]
  reg [63:0] mstatus; // @[CSR.scala 27:26]
  reg [63:0] mepc; // @[CSR.scala 28:26]
  reg [63:0] mcycle; // @[CSR.scala 29:26]
  reg [63:0] mie; // @[CSR.scala 31:26]
  reg [63:0] mscratch; // @[CSR.scala 33:26]
  wire [63:0] _mcycle_T_1 = mcycle + 64'h1; // @[CSR.scala 92:20]
  reg  intr_state; // @[CSR.scala 101:27]
  reg  mtip; // @[CSR.scala 106:21]
  reg  valid_REG; // @[CSR.scala 110:37]
  reg  valid_REG_1; // @[CSR.scala 110:60]
  wire  valid = io_mem_en ? valid_REG : valid_REG_1; // @[CSR.scala 110:18]
  wire  intr_global_en = mstatus[3]; // @[CSR.scala 115:32]
  wire  intr_clint_en = mie[7] & mtip; // @[CSR.scala 116:39]
  wire  _T = ~intr_state; // @[Conditional.scala 37:30]
  wire  _GEN_0 = intr_global_en & intr_clint_en | intr_state; // @[CSR.scala 119:46 CSR.scala 120:20 CSR.scala 101:27]
  wire [50:0] mstatus_hi_hi_hi = mstatus[63:13]; // @[CSR.scala 129:31]
  wire [2:0] mstatus_hi_lo_lo = mstatus[10:8]; // @[CSR.scala 129:58]
  wire [2:0] mstatus_lo_hi_lo = mstatus[6:4]; // @[CSR.scala 129:86]
  wire [2:0] mstatus_lo_lo_lo = mstatus[2:0]; // @[CSR.scala 129:106]
  wire [63:0] _mstatus_T = {mstatus_hi_hi_hi,1'h1,1'h1,mstatus_hi_lo_lo,intr_global_en,mstatus_lo_hi_lo,1'h0,
    mstatus_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_2 = valid ? {{32'd0}, io_pc} : mepc; // @[CSR.scala 125:20 CSR.scala 127:14 CSR.scala 28:26]
  wire [63:0] _GEN_3 = valid ? 64'h8000000000000007 : mcause; // @[CSR.scala 125:20 CSR.scala 128:16 CSR.scala 26:26]
  wire [63:0] _GEN_4 = valid ? _mstatus_T : mstatus; // @[CSR.scala 125:20 CSR.scala 129:17 CSR.scala 27:26]
  wire [63:0] _GEN_8 = intr_state ? _GEN_2 : mepc; // @[Conditional.scala 39:67 CSR.scala 28:26]
  wire [63:0] _GEN_9 = intr_state ? _GEN_3 : mcause; // @[Conditional.scala 39:67 CSR.scala 26:26]
  wire [63:0] _GEN_10 = intr_state ? _GEN_4 : mstatus; // @[Conditional.scala 39:67 CSR.scala 27:26]
  wire [63:0] _GEN_16 = _T ? mepc : _GEN_8; // @[Conditional.scala 40:58 CSR.scala 28:26]
  wire [63:0] _GEN_17 = _T ? mcause : _GEN_9; // @[Conditional.scala 40:58 CSR.scala 26:26]
  wire [63:0] _GEN_18 = _T ? mstatus : _GEN_10; // @[Conditional.scala 40:58 CSR.scala 27:26]
  wire  _io_csr_data_T = io_fuType == 3'h3; // @[CSR.scala 138:36]
  wire  _io_csr_data_T_2 = io_fuType == 3'h3 & ~io_irq; // @[CSR.scala 138:47]
  wire [63:0] _io_csr_data_rdata_T_1 = 12'h305 == io_rs2[11:0] ? mtvec : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_csr_data_rdata_T_3 = 12'h342 == io_rs2[11:0] ? mcause : _io_csr_data_rdata_T_1; // @[Mux.scala 80:57]
  wire [63:0] _io_csr_data_rdata_T_5 = 12'h341 == io_rs2[11:0] ? mepc : _io_csr_data_rdata_T_3; // @[Mux.scala 80:57]
  wire [63:0] _io_csr_data_rdata_T_7 = 12'h300 == io_rs2[11:0] ? mstatus : _io_csr_data_rdata_T_5; // @[Mux.scala 80:57]
  wire [63:0] _io_csr_data_rdata_T_9 = 12'hb00 == io_rs2[11:0] ? mcycle : _io_csr_data_rdata_T_7; // @[Mux.scala 80:57]
  wire [63:0] _io_csr_data_rdata_T_11 = 12'hb02 == io_rs2[11:0] ? 64'h0 : _io_csr_data_rdata_T_9; // @[Mux.scala 80:57]
  wire [63:0] _io_csr_data_rdata_T_13 = 12'h340 == io_rs2[11:0] ? mscratch : _io_csr_data_rdata_T_11; // @[Mux.scala 80:57]
  wire [63:0] io_csr_data_rdata = 12'h304 == io_rs2[11:0] ? mie : _io_csr_data_rdata_T_13; // @[Mux.scala 80:57]
  wire [63:0] _io_csr_data_wdata_T = io_csr_data_rdata | io_rs1; // @[CSR.scala 48:23]
  wire [63:0] _io_csr_data_wdata_T_1 = ~io_rs1; // @[CSR.scala 49:25]
  wire [63:0] _io_csr_data_wdata_T_2 = io_csr_data_rdata & _io_csr_data_wdata_T_1; // @[CSR.scala 49:23]
  wire [63:0] _io_csr_data_wdata_T_7 = 6'h2c == io_op_type ? io_rs1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_csr_data_wdata_T_9 = 6'h2d == io_op_type ? _io_csr_data_wdata_T : _io_csr_data_wdata_T_7; // @[Mux.scala 80:57]
  wire [63:0] _io_csr_data_wdata_T_11 = 6'h2e == io_op_type ? _io_csr_data_wdata_T_2 : _io_csr_data_wdata_T_9; // @[Mux.scala 80:57]
  wire [63:0] _io_csr_data_wdata_T_13 = 6'h2f == io_op_type ? io_rs1 : _io_csr_data_wdata_T_11; // @[Mux.scala 80:57]
  wire [63:0] _io_csr_data_wdata_T_15 = 6'h30 == io_op_type ? _io_csr_data_wdata_T : _io_csr_data_wdata_T_13; // @[Mux.scala 80:57]
  wire [63:0] io_csr_data_wdata = 6'h31 == io_op_type ? _io_csr_data_wdata_T_2 : _io_csr_data_wdata_T_15; // @[Mux.scala 80:57]
  wire [1:0] io_csr_data_mstatus_xs = io_csr_data_wdata[16:15]; // @[CSR.scala 58:31]
  wire [1:0] io_csr_data_mstatus_fs = io_csr_data_wdata[14:13]; // @[CSR.scala 59:31]
  wire  io_csr_data_mstatus_hi = io_csr_data_mstatus_xs == 2'h3 | io_csr_data_mstatus_fs == 2'h3; // @[CSR.scala 60:52]
  wire [62:0] io_csr_data_mstatus_lo = io_csr_data_wdata[62:0]; // @[CSR.scala 61:41]
  wire [63:0] _io_csr_data_mstatus_T = {io_csr_data_mstatus_hi,io_csr_data_mstatus_lo}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_22 = io_rs2[11:0] == 12'h300 ? _io_csr_data_mstatus_T : _GEN_18; // @[CSR.scala 57:33 CSR.scala 61:17]
  wire  io_csr_Jmp_en_br_en = _io_csr_data_T & io_op_type == 6'h32; // @[CSR.scala 72:23]
  wire  io_csr_Jmp_en_mstatus_lo_lo_hi = mstatus[7]; // @[CSR.scala 78:92]
  wire [63:0] _io_csr_Jmp_en_mstatus_T_1 = {mstatus_hi_hi_hi,1'h0,1'h0,mstatus_hi_lo_lo,1'h1,mstatus_lo_hi_lo,
    io_csr_Jmp_en_mstatus_lo_lo_hi,mstatus_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] _io_csr_Jmp_addr_br_addr_T_1 = 12'h0 == io_rs2[11:0] ? mtvec : 64'h80000000; // @[Mux.scala 80:57]
  wire [63:0] io_csr_Jmp_addr_br_addr = 12'h302 == io_rs2[11:0] ? mepc : _io_csr_Jmp_addr_br_addr_T_1; // @[Mux.scala 80:57]
  wire [63:0] _io_csr_Jmp_addr_T_1 = io_irq ? mtvec : io_csr_Jmp_addr_br_addr; // @[CSR.scala 140:25]
  assign io_csr_Jmp_addr = _io_csr_Jmp_addr_T_1[31:0]; // @[CSR.scala 140:19]
  assign io_csr_Jmp_en = io_csr_Jmp_en_br_en | io_irq; // @[CSR.scala 139:84]
  assign io_csr_data = 12'h304 == io_rs2[11:0] ? mie : _io_csr_data_rdata_T_13; // @[Mux.scala 80:57]
  assign io_irq = intr_state & valid; // @[CSR.scala 137:37]
  always @(posedge clock) begin
    if (reset) begin // @[CSR.scala 25:26]
      mtvec <= 64'h0; // @[CSR.scala 25:26]
    end else if (_io_csr_data_T_2 & io_op_type != 6'h32) begin // @[CSR.scala 55:36]
      if (io_rs2[11:0] == 12'h305) begin // @[CSR.scala 56:31]
        if (6'h31 == io_op_type) begin // @[Mux.scala 80:57]
          mtvec <= _io_csr_data_wdata_T_2;
        end else begin
          mtvec <= _io_csr_data_wdata_T_15;
        end
      end
    end
    if (reset) begin // @[CSR.scala 26:26]
      mcause <= 64'h0; // @[CSR.scala 26:26]
    end else if (io_csr_Jmp_en_br_en & io_rs2[11:0] == 12'h0) begin // @[CSR.scala 73:40]
      mcause <= 64'hb; // @[CSR.scala 75:14]
    end else if (_io_csr_data_T_2 & io_op_type != 6'h32) begin // @[CSR.scala 55:36]
      if (io_rs2[11:0] == 12'h342) begin // @[CSR.scala 63:32]
        mcause <= io_csr_data_wdata; // @[CSR.scala 63:41]
      end else begin
        mcause <= _GEN_17;
      end
    end else begin
      mcause <= _GEN_17;
    end
    if (reset) begin // @[CSR.scala 27:26]
      mstatus <= 64'h1800; // @[CSR.scala 27:26]
    end else if (io_csr_Jmp_en_br_en & io_rs2[11:0] == 12'h0) begin // @[CSR.scala 73:40]
      mstatus <= _mstatus_T; // @[CSR.scala 76:15]
    end else if (io_csr_Jmp_en_br_en & io_rs2[11:0] == 12'h302) begin // @[CSR.scala 77:45]
      mstatus <= _io_csr_Jmp_en_mstatus_T_1; // @[CSR.scala 78:15]
    end else if (_io_csr_data_T_2 & io_op_type != 6'h32) begin // @[CSR.scala 55:36]
      mstatus <= _GEN_22;
    end else begin
      mstatus <= _GEN_18;
    end
    if (reset) begin // @[CSR.scala 28:26]
      mepc <= 64'h0; // @[CSR.scala 28:26]
    end else if (io_csr_Jmp_en_br_en & io_rs2[11:0] == 12'h0) begin // @[CSR.scala 73:40]
      mepc <= {{32'd0}, io_pc}; // @[CSR.scala 74:12]
    end else if (_io_csr_data_T_2 & io_op_type != 6'h32) begin // @[CSR.scala 55:36]
      if (io_rs2[11:0] == 12'h341) begin // @[CSR.scala 62:30]
        mepc <= io_csr_data_wdata; // @[CSR.scala 62:37]
      end else begin
        mepc <= _GEN_16;
      end
    end else begin
      mepc <= _GEN_16;
    end
    if (reset) begin // @[CSR.scala 29:26]
      mcycle <= 64'h0; // @[CSR.scala 29:26]
    end else begin
      mcycle <= _mcycle_T_1; // @[CSR.scala 92:10]
    end
    if (reset) begin // @[CSR.scala 31:26]
      mie <= 64'h0; // @[CSR.scala 31:26]
    end else if (_io_csr_data_T_2 & io_op_type != 6'h32) begin // @[CSR.scala 55:36]
      if (io_rs2[11:0] == 12'h304) begin // @[CSR.scala 64:29]
        if (6'h31 == io_op_type) begin // @[Mux.scala 80:57]
          mie <= _io_csr_data_wdata_T_2;
        end else begin
          mie <= _io_csr_data_wdata_T_15;
        end
      end
    end
    if (reset) begin // @[CSR.scala 33:26]
      mscratch <= 64'h0; // @[CSR.scala 33:26]
    end else if (_io_csr_data_T_2 & io_op_type != 6'h32) begin // @[CSR.scala 55:36]
      if (io_rs2[11:0] == 12'h340) begin // @[CSR.scala 65:34]
        if (6'h31 == io_op_type) begin // @[Mux.scala 80:57]
          mscratch <= _io_csr_data_wdata_T_2;
        end else begin
          mscratch <= _io_csr_data_wdata_T_15;
        end
      end
    end
    if (reset) begin // @[CSR.scala 101:27]
      intr_state <= 1'h0; // @[CSR.scala 101:27]
    end else if (_T) begin // @[Conditional.scala 40:58]
      intr_state <= _GEN_0;
    end else if (intr_state) begin // @[Conditional.scala 39:67]
      if (valid) begin // @[CSR.scala 125:20]
        intr_state <= 1'h0; // @[CSR.scala 132:20]
      end
    end
    if (reset) begin // @[CSR.scala 106:21]
      mtip <= 1'h0; // @[CSR.scala 106:21]
    end else begin
      mtip <= mtip_0;
    end
    valid_REG <= io_mem_valid; // @[CSR.scala 110:37]
    valid_REG_1 <= io_if_valid; // @[CSR.scala 110:60]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtvec = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mcause = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mstatus = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mepc = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mcycle = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mie = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mscratch = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  intr_state = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  mtip = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  valid_REG = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  valid_REG_1 = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210340_Cache_1(
  input         clock,
  input         reset,
  output [5:0]   io_sram4_addr,
  output         io_sram4_cen,
  output         io_sram4_wen,
  output [127:0] io_sram4_wdata,
  input  [127:0] io_sram4_rdata,
  output [5:0]   io_sram5_addr,
  output         io_sram5_cen,
  output         io_sram5_wen,
  output [127:0] io_sram5_wdata,
  input  [127:0] io_sram5_rdata,
  output [5:0]   io_sram6_addr,
  output         io_sram6_cen,
  output         io_sram6_wen,
  output [127:0] io_sram6_wdata,
  input  [127:0] io_sram6_rdata,
  output [5:0]   io_sram7_addr,
  output         io_sram7_cen,
  output         io_sram7_wen,
  output [127:0] io_sram7_wdata,
  input  [127:0] io_sram7_rdata,  
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output        io_out_req_bits_aen,
  output        io_out_req_bits_ren,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_req_bits_wlast,
  output        io_out_req_bits_wen,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata,
  input         io_out_resp_bits_rlast,
  input         fence_i_0,
  output        dcache_fi_complete_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [127:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [127:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [63:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [127:0] _RAND_213;
  reg [31:0] _RAND_214;
`endif // RANDOMIZE_REG_INIT
  // wire  sram_0_clock; // @[Cache.scala 91:22]
  wire  sram_0_io_en; // @[Cache.scala 91:22]
  wire  sram_0_io_wen; // @[Cache.scala 91:22]
  wire [5:0] sram_0_io_addr; // @[Cache.scala 91:22]
  wire [127:0] sram_0_io_wdata; // @[Cache.scala 91:22]
  wire [127:0] sram_0_io_rdata; // @[Cache.scala 91:22]
  // wire  sram_1_clock; // @[Cache.scala 91:22]
  wire  sram_1_io_en; // @[Cache.scala 91:22]
  wire  sram_1_io_wen; // @[Cache.scala 91:22]
  wire [5:0] sram_1_io_addr; // @[Cache.scala 91:22]
  wire [127:0] sram_1_io_wdata; // @[Cache.scala 91:22]
  wire [127:0] sram_1_io_rdata; // @[Cache.scala 91:22]
  // wire  sram_2_clock; // @[Cache.scala 91:22]
  wire  sram_2_io_en; // @[Cache.scala 91:22]
  wire  sram_2_io_wen; // @[Cache.scala 91:22]
  wire [5:0] sram_2_io_addr; // @[Cache.scala 91:22]
  wire [127:0] sram_2_io_wdata; // @[Cache.scala 91:22]
  wire [127:0] sram_2_io_rdata; // @[Cache.scala 91:22]
  // wire  sram_3_clock; // @[Cache.scala 91:22]
  wire  sram_3_io_en; // @[Cache.scala 91:22]
  wire  sram_3_io_wen; // @[Cache.scala 91:22]
  wire [5:0] sram_3_io_addr; // @[Cache.scala 91:22]
  wire [127:0] sram_3_io_wdata; // @[Cache.scala 91:22]
  wire [127:0] sram_3_io_rdata; // @[Cache.scala 91:22]
  wire  meta_0_clock; // @[Cache.scala 99:22]
  wire  meta_0_reset; // @[Cache.scala 99:22]
  wire [5:0] meta_0_io_idx; // @[Cache.scala 99:22]
  wire [20:0] meta_0_io_tag_r; // @[Cache.scala 99:22]
  wire [20:0] meta_0_io_tag_w; // @[Cache.scala 99:22]
  wire  meta_0_io_tag_wen; // @[Cache.scala 99:22]
  wire  meta_0_io_dirty_r; // @[Cache.scala 99:22]
  wire  meta_0_io_dirty_w; // @[Cache.scala 99:22]
  wire  meta_0_io_dirty_wen; // @[Cache.scala 99:22]
  wire  meta_0_io_valid_r; // @[Cache.scala 99:22]
  wire  meta_0_io_invalidate; // @[Cache.scala 99:22]
  wire  meta_0_io_dirty_r_async; // @[Cache.scala 99:22]
  wire  meta_0_io_valid_r_async; // @[Cache.scala 99:22]
  wire  meta_1_clock; // @[Cache.scala 99:22]
  wire  meta_1_reset; // @[Cache.scala 99:22]
  wire [5:0] meta_1_io_idx; // @[Cache.scala 99:22]
  wire [20:0] meta_1_io_tag_r; // @[Cache.scala 99:22]
  wire [20:0] meta_1_io_tag_w; // @[Cache.scala 99:22]
  wire  meta_1_io_tag_wen; // @[Cache.scala 99:22]
  wire  meta_1_io_dirty_r; // @[Cache.scala 99:22]
  wire  meta_1_io_dirty_w; // @[Cache.scala 99:22]
  wire  meta_1_io_dirty_wen; // @[Cache.scala 99:22]
  wire  meta_1_io_valid_r; // @[Cache.scala 99:22]
  wire  meta_1_io_invalidate; // @[Cache.scala 99:22]
  wire  meta_1_io_dirty_r_async; // @[Cache.scala 99:22]
  wire  meta_1_io_valid_r_async; // @[Cache.scala 99:22]
  wire  meta_2_clock; // @[Cache.scala 99:22]
  wire  meta_2_reset; // @[Cache.scala 99:22]
  wire [5:0] meta_2_io_idx; // @[Cache.scala 99:22]
  wire [20:0] meta_2_io_tag_r; // @[Cache.scala 99:22]
  wire [20:0] meta_2_io_tag_w; // @[Cache.scala 99:22]
  wire  meta_2_io_tag_wen; // @[Cache.scala 99:22]
  wire  meta_2_io_dirty_r; // @[Cache.scala 99:22]
  wire  meta_2_io_dirty_w; // @[Cache.scala 99:22]
  wire  meta_2_io_dirty_wen; // @[Cache.scala 99:22]
  wire  meta_2_io_valid_r; // @[Cache.scala 99:22]
  wire  meta_2_io_invalidate; // @[Cache.scala 99:22]
  wire  meta_2_io_dirty_r_async; // @[Cache.scala 99:22]
  wire  meta_2_io_valid_r_async; // @[Cache.scala 99:22]
  wire  meta_3_clock; // @[Cache.scala 99:22]
  wire  meta_3_reset; // @[Cache.scala 99:22]
  wire [5:0] meta_3_io_idx; // @[Cache.scala 99:22]
  wire [20:0] meta_3_io_tag_r; // @[Cache.scala 99:22]
  wire [20:0] meta_3_io_tag_w; // @[Cache.scala 99:22]
  wire  meta_3_io_tag_wen; // @[Cache.scala 99:22]
  wire  meta_3_io_dirty_r; // @[Cache.scala 99:22]
  wire  meta_3_io_dirty_w; // @[Cache.scala 99:22]
  wire  meta_3_io_dirty_wen; // @[Cache.scala 99:22]
  wire  meta_3_io_valid_r; // @[Cache.scala 99:22]
  wire  meta_3_io_invalidate; // @[Cache.scala 99:22]
  wire  meta_3_io_dirty_r_async; // @[Cache.scala 99:22]
  wire  meta_3_io_valid_r_async; // @[Cache.scala 99:22]
  reg  plru0_0; // @[Cache.scala 131:22]
  reg  plru0_1; // @[Cache.scala 131:22]
  reg  plru0_2; // @[Cache.scala 131:22]
  reg  plru0_3; // @[Cache.scala 131:22]
  reg  plru0_4; // @[Cache.scala 131:22]
  reg  plru0_5; // @[Cache.scala 131:22]
  reg  plru0_6; // @[Cache.scala 131:22]
  reg  plru0_7; // @[Cache.scala 131:22]
  reg  plru0_8; // @[Cache.scala 131:22]
  reg  plru0_9; // @[Cache.scala 131:22]
  reg  plru0_10; // @[Cache.scala 131:22]
  reg  plru0_11; // @[Cache.scala 131:22]
  reg  plru0_12; // @[Cache.scala 131:22]
  reg  plru0_13; // @[Cache.scala 131:22]
  reg  plru0_14; // @[Cache.scala 131:22]
  reg  plru0_15; // @[Cache.scala 131:22]
  reg  plru0_16; // @[Cache.scala 131:22]
  reg  plru0_17; // @[Cache.scala 131:22]
  reg  plru0_18; // @[Cache.scala 131:22]
  reg  plru0_19; // @[Cache.scala 131:22]
  reg  plru0_20; // @[Cache.scala 131:22]
  reg  plru0_21; // @[Cache.scala 131:22]
  reg  plru0_22; // @[Cache.scala 131:22]
  reg  plru0_23; // @[Cache.scala 131:22]
  reg  plru0_24; // @[Cache.scala 131:22]
  reg  plru0_25; // @[Cache.scala 131:22]
  reg  plru0_26; // @[Cache.scala 131:22]
  reg  plru0_27; // @[Cache.scala 131:22]
  reg  plru0_28; // @[Cache.scala 131:22]
  reg  plru0_29; // @[Cache.scala 131:22]
  reg  plru0_30; // @[Cache.scala 131:22]
  reg  plru0_31; // @[Cache.scala 131:22]
  reg  plru0_32; // @[Cache.scala 131:22]
  reg  plru0_33; // @[Cache.scala 131:22]
  reg  plru0_34; // @[Cache.scala 131:22]
  reg  plru0_35; // @[Cache.scala 131:22]
  reg  plru0_36; // @[Cache.scala 131:22]
  reg  plru0_37; // @[Cache.scala 131:22]
  reg  plru0_38; // @[Cache.scala 131:22]
  reg  plru0_39; // @[Cache.scala 131:22]
  reg  plru0_40; // @[Cache.scala 131:22]
  reg  plru0_41; // @[Cache.scala 131:22]
  reg  plru0_42; // @[Cache.scala 131:22]
  reg  plru0_43; // @[Cache.scala 131:22]
  reg  plru0_44; // @[Cache.scala 131:22]
  reg  plru0_45; // @[Cache.scala 131:22]
  reg  plru0_46; // @[Cache.scala 131:22]
  reg  plru0_47; // @[Cache.scala 131:22]
  reg  plru0_48; // @[Cache.scala 131:22]
  reg  plru0_49; // @[Cache.scala 131:22]
  reg  plru0_50; // @[Cache.scala 131:22]
  reg  plru0_51; // @[Cache.scala 131:22]
  reg  plru0_52; // @[Cache.scala 131:22]
  reg  plru0_53; // @[Cache.scala 131:22]
  reg  plru0_54; // @[Cache.scala 131:22]
  reg  plru0_55; // @[Cache.scala 131:22]
  reg  plru0_56; // @[Cache.scala 131:22]
  reg  plru0_57; // @[Cache.scala 131:22]
  reg  plru0_58; // @[Cache.scala 131:22]
  reg  plru0_59; // @[Cache.scala 131:22]
  reg  plru0_60; // @[Cache.scala 131:22]
  reg  plru0_61; // @[Cache.scala 131:22]
  reg  plru0_62; // @[Cache.scala 131:22]
  reg  plru0_63; // @[Cache.scala 131:22]
  reg  plru1_0; // @[Cache.scala 133:22]
  reg  plru1_1; // @[Cache.scala 133:22]
  reg  plru1_2; // @[Cache.scala 133:22]
  reg  plru1_3; // @[Cache.scala 133:22]
  reg  plru1_4; // @[Cache.scala 133:22]
  reg  plru1_5; // @[Cache.scala 133:22]
  reg  plru1_6; // @[Cache.scala 133:22]
  reg  plru1_7; // @[Cache.scala 133:22]
  reg  plru1_8; // @[Cache.scala 133:22]
  reg  plru1_9; // @[Cache.scala 133:22]
  reg  plru1_10; // @[Cache.scala 133:22]
  reg  plru1_11; // @[Cache.scala 133:22]
  reg  plru1_12; // @[Cache.scala 133:22]
  reg  plru1_13; // @[Cache.scala 133:22]
  reg  plru1_14; // @[Cache.scala 133:22]
  reg  plru1_15; // @[Cache.scala 133:22]
  reg  plru1_16; // @[Cache.scala 133:22]
  reg  plru1_17; // @[Cache.scala 133:22]
  reg  plru1_18; // @[Cache.scala 133:22]
  reg  plru1_19; // @[Cache.scala 133:22]
  reg  plru1_20; // @[Cache.scala 133:22]
  reg  plru1_21; // @[Cache.scala 133:22]
  reg  plru1_22; // @[Cache.scala 133:22]
  reg  plru1_23; // @[Cache.scala 133:22]
  reg  plru1_24; // @[Cache.scala 133:22]
  reg  plru1_25; // @[Cache.scala 133:22]
  reg  plru1_26; // @[Cache.scala 133:22]
  reg  plru1_27; // @[Cache.scala 133:22]
  reg  plru1_28; // @[Cache.scala 133:22]
  reg  plru1_29; // @[Cache.scala 133:22]
  reg  plru1_30; // @[Cache.scala 133:22]
  reg  plru1_31; // @[Cache.scala 133:22]
  reg  plru1_32; // @[Cache.scala 133:22]
  reg  plru1_33; // @[Cache.scala 133:22]
  reg  plru1_34; // @[Cache.scala 133:22]
  reg  plru1_35; // @[Cache.scala 133:22]
  reg  plru1_36; // @[Cache.scala 133:22]
  reg  plru1_37; // @[Cache.scala 133:22]
  reg  plru1_38; // @[Cache.scala 133:22]
  reg  plru1_39; // @[Cache.scala 133:22]
  reg  plru1_40; // @[Cache.scala 133:22]
  reg  plru1_41; // @[Cache.scala 133:22]
  reg  plru1_42; // @[Cache.scala 133:22]
  reg  plru1_43; // @[Cache.scala 133:22]
  reg  plru1_44; // @[Cache.scala 133:22]
  reg  plru1_45; // @[Cache.scala 133:22]
  reg  plru1_46; // @[Cache.scala 133:22]
  reg  plru1_47; // @[Cache.scala 133:22]
  reg  plru1_48; // @[Cache.scala 133:22]
  reg  plru1_49; // @[Cache.scala 133:22]
  reg  plru1_50; // @[Cache.scala 133:22]
  reg  plru1_51; // @[Cache.scala 133:22]
  reg  plru1_52; // @[Cache.scala 133:22]
  reg  plru1_53; // @[Cache.scala 133:22]
  reg  plru1_54; // @[Cache.scala 133:22]
  reg  plru1_55; // @[Cache.scala 133:22]
  reg  plru1_56; // @[Cache.scala 133:22]
  reg  plru1_57; // @[Cache.scala 133:22]
  reg  plru1_58; // @[Cache.scala 133:22]
  reg  plru1_59; // @[Cache.scala 133:22]
  reg  plru1_60; // @[Cache.scala 133:22]
  reg  plru1_61; // @[Cache.scala 133:22]
  reg  plru1_62; // @[Cache.scala 133:22]
  reg  plru1_63; // @[Cache.scala 133:22]
  reg  plru2_0; // @[Cache.scala 135:22]
  reg  plru2_1; // @[Cache.scala 135:22]
  reg  plru2_2; // @[Cache.scala 135:22]
  reg  plru2_3; // @[Cache.scala 135:22]
  reg  plru2_4; // @[Cache.scala 135:22]
  reg  plru2_5; // @[Cache.scala 135:22]
  reg  plru2_6; // @[Cache.scala 135:22]
  reg  plru2_7; // @[Cache.scala 135:22]
  reg  plru2_8; // @[Cache.scala 135:22]
  reg  plru2_9; // @[Cache.scala 135:22]
  reg  plru2_10; // @[Cache.scala 135:22]
  reg  plru2_11; // @[Cache.scala 135:22]
  reg  plru2_12; // @[Cache.scala 135:22]
  reg  plru2_13; // @[Cache.scala 135:22]
  reg  plru2_14; // @[Cache.scala 135:22]
  reg  plru2_15; // @[Cache.scala 135:22]
  reg  plru2_16; // @[Cache.scala 135:22]
  reg  plru2_17; // @[Cache.scala 135:22]
  reg  plru2_18; // @[Cache.scala 135:22]
  reg  plru2_19; // @[Cache.scala 135:22]
  reg  plru2_20; // @[Cache.scala 135:22]
  reg  plru2_21; // @[Cache.scala 135:22]
  reg  plru2_22; // @[Cache.scala 135:22]
  reg  plru2_23; // @[Cache.scala 135:22]
  reg  plru2_24; // @[Cache.scala 135:22]
  reg  plru2_25; // @[Cache.scala 135:22]
  reg  plru2_26; // @[Cache.scala 135:22]
  reg  plru2_27; // @[Cache.scala 135:22]
  reg  plru2_28; // @[Cache.scala 135:22]
  reg  plru2_29; // @[Cache.scala 135:22]
  reg  plru2_30; // @[Cache.scala 135:22]
  reg  plru2_31; // @[Cache.scala 135:22]
  reg  plru2_32; // @[Cache.scala 135:22]
  reg  plru2_33; // @[Cache.scala 135:22]
  reg  plru2_34; // @[Cache.scala 135:22]
  reg  plru2_35; // @[Cache.scala 135:22]
  reg  plru2_36; // @[Cache.scala 135:22]
  reg  plru2_37; // @[Cache.scala 135:22]
  reg  plru2_38; // @[Cache.scala 135:22]
  reg  plru2_39; // @[Cache.scala 135:22]
  reg  plru2_40; // @[Cache.scala 135:22]
  reg  plru2_41; // @[Cache.scala 135:22]
  reg  plru2_42; // @[Cache.scala 135:22]
  reg  plru2_43; // @[Cache.scala 135:22]
  reg  plru2_44; // @[Cache.scala 135:22]
  reg  plru2_45; // @[Cache.scala 135:22]
  reg  plru2_46; // @[Cache.scala 135:22]
  reg  plru2_47; // @[Cache.scala 135:22]
  reg  plru2_48; // @[Cache.scala 135:22]
  reg  plru2_49; // @[Cache.scala 135:22]
  reg  plru2_50; // @[Cache.scala 135:22]
  reg  plru2_51; // @[Cache.scala 135:22]
  reg  plru2_52; // @[Cache.scala 135:22]
  reg  plru2_53; // @[Cache.scala 135:22]
  reg  plru2_54; // @[Cache.scala 135:22]
  reg  plru2_55; // @[Cache.scala 135:22]
  reg  plru2_56; // @[Cache.scala 135:22]
  reg  plru2_57; // @[Cache.scala 135:22]
  reg  plru2_58; // @[Cache.scala 135:22]
  reg  plru2_59; // @[Cache.scala 135:22]
  reg  plru2_60; // @[Cache.scala 135:22]
  reg  plru2_61; // @[Cache.scala 135:22]
  reg  plru2_62; // @[Cache.scala 135:22]
  reg  plru2_63; // @[Cache.scala 135:22]
  reg  s2_hit_real_REG; // @[Cache.scala 263:32]
  wire [20:0] tag_out_0 = meta_0_io_tag_r;
  reg [31:0] s2_addr; // @[Cache.scala 209:25]
  wire [20:0] s2_tag = s2_addr[30:10]; // @[Cache.scala 212:25]
  wire  valid_out_0 = meta_0_io_valid_r;
  wire  hit_0 = tag_out_0 == s2_tag & valid_out_0; // @[Cache.scala 222:25]
  wire [20:0] tag_out_1 = meta_1_io_tag_r;
  wire  valid_out_1 = meta_1_io_valid_r;
  wire  hit_1 = tag_out_1 == s2_tag & valid_out_1; // @[Cache.scala 222:25]
  wire [20:0] tag_out_2 = meta_2_io_tag_r;
  wire  valid_out_2 = meta_2_io_valid_r;
  wire  hit_2 = tag_out_2 == s2_tag & valid_out_2; // @[Cache.scala 222:25]
  wire [20:0] tag_out_3 = meta_3_io_tag_r;
  wire  valid_out_3 = meta_3_io_valid_r;
  wire  hit_3 = tag_out_3 == s2_tag & valid_out_3; // @[Cache.scala 222:25]
  wire [3:0] _s2_hit_T = {hit_0,hit_1,hit_2,hit_3}; // @[Cat.scala 30:58]
  wire  s2_hit = |_s2_hit_T; // @[Cache.scala 224:25]
  reg  s2_reg_hit; // @[Cache.scala 231:27]
  wire  s2_hit_real = s2_hit_real_REG ? s2_hit : s2_reg_hit; // @[Cache.scala 263:24]
  reg  s2_wen; // @[Cache.scala 213:25]
  reg [3:0] state; // @[Cache.scala 207:22]
  wire  _hit_ready_T = state == 4'h7; // @[Cache.scala 265:37]
  wire  _hit_ready_T_2 = s2_wen ? state == 4'h7 : state == 4'h0; // @[Cache.scala 265:22]
  wire  hit_ready = s2_hit_real & _hit_ready_T_2; // @[Cache.scala 264:31]
  wire  invalid_ready = state == 4'h8; // @[Cache.scala 267:30]
  wire  fi_ready = (hit_ready | _hit_ready_T) & io_in_resp_ready | invalid_ready; // @[Cache.scala 270:66]
  reg  fi_valid; // @[ID.scala 18:20]
  wire  _GEN_0 = fence_i_0 | fi_valid; // @[ID.scala 24:20 ID.scala 24:24 ID.scala 18:20]
  reg [2:0] fi_state; // @[Cache.scala 399:25]
  wire  _T_34 = 3'h0 == fi_state; // @[Conditional.scala 37:30]
  wire  _T_35 = 3'h1 == fi_state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h2 == fi_state; // @[Conditional.scala 37:30]
  wire  _T_43 = 3'h3 == fi_state; // @[Conditional.scala 37:30]
  wire  _T_45 = 3'h4 == fi_state; // @[Conditional.scala 37:30]
  wire  _T_48 = 3'h5 == fi_state; // @[Conditional.scala 37:30]
  wire  _GEN_3563 = _T_45 ? 1'h0 : _T_48; // @[Conditional.scala 39:67]
  wire  _GEN_3566 = _T_43 ? 1'h0 : _GEN_3563; // @[Conditional.scala 39:67]
  wire  _GEN_3569 = _T_41 ? 1'h0 : _GEN_3566; // @[Conditional.scala 39:67]
  wire  _GEN_3576 = _T_35 ? 1'h0 : _GEN_3569; // @[Conditional.scala 39:67]
  wire  dcache_fi_complete = _T_34 ? 1'h0 : _GEN_3576; // @[Conditional.scala 40:58]
  wire  fi_fire = fi_valid & fi_ready; // @[Cache.scala 163:26]
  wire [5:0] s1_idx = io_in_req_bits_addr[9:4]; // @[Cache.scala 171:25]
  wire [5:0] _GEN_3 = fi_ready ? s1_idx : 6'h0; // @[Cache.scala 181:24 Cache.scala 184:17 Cache.scala 111:15]
  wire  s2_offs = s2_addr[3]; // @[Cache.scala 210:25]
  wire [5:0] s2_idx = s2_addr[9:4]; // @[Cache.scala 211:25]
  reg [63:0] s2_wdata; // @[Cache.scala 214:25]
  reg [7:0] s2_wmask; // @[Cache.scala 215:25]
  wire [3:0] _s2_way_T = {hit_3,hit_2,hit_1,hit_0}; // @[OneHot.scala 22:45]
  wire [1:0] s2_way_hi_1 = _s2_way_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] s2_way_lo_1 = _s2_way_T[1:0]; // @[OneHot.scala 31:18]
  wire  s2_way_hi_2 = |s2_way_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _s2_way_T_1 = s2_way_hi_1 | s2_way_lo_1; // @[OneHot.scala 32:28]
  wire  s2_way_lo_2 = _s2_way_T_1[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] s2_way = {s2_way_hi_2,s2_way_lo_2}; // @[Cat.scala 30:58]
  reg [127:0] s2_reg_rdata; // @[Cache.scala 233:29]
  reg  s2_reg_dirty; // @[Cache.scala 234:29]
  reg [20:0] s2_reg_tag_r; // @[Cache.scala 235:29]
  reg [127:0] s2_reg_dat_w; // @[Cache.scala 236:29]
  reg  REG; // @[Cache.scala 244:41]
  wire [127:0] sram_out_0 = sram_0_io_rdata;
  wire [127:0] sram_out_1 = sram_1_io_rdata;
  wire [127:0] _GEN_5 = 2'h1 == s2_way ? sram_out_1 : sram_out_0; // @[Cache.scala 249:18 Cache.scala 249:18]
  wire [127:0] sram_out_2 = sram_2_io_rdata;
  wire [127:0] _GEN_6 = 2'h2 == s2_way ? sram_out_2 : _GEN_5; // @[Cache.scala 249:18 Cache.scala 249:18]
  wire [127:0] sram_out_3 = sram_3_io_rdata;
  wire [127:0] _GEN_7 = 2'h3 == s2_way ? sram_out_3 : _GEN_6; // @[Cache.scala 249:18 Cache.scala 249:18]
  wire  _GEN_37 = 6'h1 == s2_idx ? plru0_1 : plru0_0; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_38 = 6'h2 == s2_idx ? plru0_2 : _GEN_37; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_39 = 6'h3 == s2_idx ? plru0_3 : _GEN_38; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_40 = 6'h4 == s2_idx ? plru0_4 : _GEN_39; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_41 = 6'h5 == s2_idx ? plru0_5 : _GEN_40; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_42 = 6'h6 == s2_idx ? plru0_6 : _GEN_41; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_43 = 6'h7 == s2_idx ? plru0_7 : _GEN_42; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_44 = 6'h8 == s2_idx ? plru0_8 : _GEN_43; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_45 = 6'h9 == s2_idx ? plru0_9 : _GEN_44; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_46 = 6'ha == s2_idx ? plru0_10 : _GEN_45; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_47 = 6'hb == s2_idx ? plru0_11 : _GEN_46; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_48 = 6'hc == s2_idx ? plru0_12 : _GEN_47; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_49 = 6'hd == s2_idx ? plru0_13 : _GEN_48; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_50 = 6'he == s2_idx ? plru0_14 : _GEN_49; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_51 = 6'hf == s2_idx ? plru0_15 : _GEN_50; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_52 = 6'h10 == s2_idx ? plru0_16 : _GEN_51; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_53 = 6'h11 == s2_idx ? plru0_17 : _GEN_52; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_54 = 6'h12 == s2_idx ? plru0_18 : _GEN_53; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_55 = 6'h13 == s2_idx ? plru0_19 : _GEN_54; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_56 = 6'h14 == s2_idx ? plru0_20 : _GEN_55; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_57 = 6'h15 == s2_idx ? plru0_21 : _GEN_56; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_58 = 6'h16 == s2_idx ? plru0_22 : _GEN_57; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_59 = 6'h17 == s2_idx ? plru0_23 : _GEN_58; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_60 = 6'h18 == s2_idx ? plru0_24 : _GEN_59; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_61 = 6'h19 == s2_idx ? plru0_25 : _GEN_60; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_62 = 6'h1a == s2_idx ? plru0_26 : _GEN_61; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_63 = 6'h1b == s2_idx ? plru0_27 : _GEN_62; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_64 = 6'h1c == s2_idx ? plru0_28 : _GEN_63; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_65 = 6'h1d == s2_idx ? plru0_29 : _GEN_64; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_66 = 6'h1e == s2_idx ? plru0_30 : _GEN_65; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_67 = 6'h1f == s2_idx ? plru0_31 : _GEN_66; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_68 = 6'h20 == s2_idx ? plru0_32 : _GEN_67; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_69 = 6'h21 == s2_idx ? plru0_33 : _GEN_68; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_70 = 6'h22 == s2_idx ? plru0_34 : _GEN_69; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_71 = 6'h23 == s2_idx ? plru0_35 : _GEN_70; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_72 = 6'h24 == s2_idx ? plru0_36 : _GEN_71; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_73 = 6'h25 == s2_idx ? plru0_37 : _GEN_72; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_74 = 6'h26 == s2_idx ? plru0_38 : _GEN_73; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_75 = 6'h27 == s2_idx ? plru0_39 : _GEN_74; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_76 = 6'h28 == s2_idx ? plru0_40 : _GEN_75; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_77 = 6'h29 == s2_idx ? plru0_41 : _GEN_76; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_78 = 6'h2a == s2_idx ? plru0_42 : _GEN_77; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_79 = 6'h2b == s2_idx ? plru0_43 : _GEN_78; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_80 = 6'h2c == s2_idx ? plru0_44 : _GEN_79; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_81 = 6'h2d == s2_idx ? plru0_45 : _GEN_80; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_82 = 6'h2e == s2_idx ? plru0_46 : _GEN_81; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_83 = 6'h2f == s2_idx ? plru0_47 : _GEN_82; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_84 = 6'h30 == s2_idx ? plru0_48 : _GEN_83; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_85 = 6'h31 == s2_idx ? plru0_49 : _GEN_84; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_86 = 6'h32 == s2_idx ? plru0_50 : _GEN_85; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_87 = 6'h33 == s2_idx ? plru0_51 : _GEN_86; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_88 = 6'h34 == s2_idx ? plru0_52 : _GEN_87; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_89 = 6'h35 == s2_idx ? plru0_53 : _GEN_88; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_90 = 6'h36 == s2_idx ? plru0_54 : _GEN_89; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_91 = 6'h37 == s2_idx ? plru0_55 : _GEN_90; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_92 = 6'h38 == s2_idx ? plru0_56 : _GEN_91; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_93 = 6'h39 == s2_idx ? plru0_57 : _GEN_92; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_94 = 6'h3a == s2_idx ? plru0_58 : _GEN_93; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_95 = 6'h3b == s2_idx ? plru0_59 : _GEN_94; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_96 = 6'h3c == s2_idx ? plru0_60 : _GEN_95; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_97 = 6'h3d == s2_idx ? plru0_61 : _GEN_96; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_98 = 6'h3e == s2_idx ? plru0_62 : _GEN_97; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_99 = 6'h3f == s2_idx ? plru0_63 : _GEN_98; // @[Cache.scala 256:40 Cache.scala 256:40]
  wire  _GEN_101 = 6'h1 == s2_idx ? plru1_1 : plru1_0; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_102 = 6'h2 == s2_idx ? plru1_2 : _GEN_101; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_103 = 6'h3 == s2_idx ? plru1_3 : _GEN_102; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_104 = 6'h4 == s2_idx ? plru1_4 : _GEN_103; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_105 = 6'h5 == s2_idx ? plru1_5 : _GEN_104; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_106 = 6'h6 == s2_idx ? plru1_6 : _GEN_105; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_107 = 6'h7 == s2_idx ? plru1_7 : _GEN_106; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_108 = 6'h8 == s2_idx ? plru1_8 : _GEN_107; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_109 = 6'h9 == s2_idx ? plru1_9 : _GEN_108; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_110 = 6'ha == s2_idx ? plru1_10 : _GEN_109; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_111 = 6'hb == s2_idx ? plru1_11 : _GEN_110; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_112 = 6'hc == s2_idx ? plru1_12 : _GEN_111; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_113 = 6'hd == s2_idx ? plru1_13 : _GEN_112; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_114 = 6'he == s2_idx ? plru1_14 : _GEN_113; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_115 = 6'hf == s2_idx ? plru1_15 : _GEN_114; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_116 = 6'h10 == s2_idx ? plru1_16 : _GEN_115; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_117 = 6'h11 == s2_idx ? plru1_17 : _GEN_116; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_118 = 6'h12 == s2_idx ? plru1_18 : _GEN_117; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_119 = 6'h13 == s2_idx ? plru1_19 : _GEN_118; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_120 = 6'h14 == s2_idx ? plru1_20 : _GEN_119; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_121 = 6'h15 == s2_idx ? plru1_21 : _GEN_120; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_122 = 6'h16 == s2_idx ? plru1_22 : _GEN_121; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_123 = 6'h17 == s2_idx ? plru1_23 : _GEN_122; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_124 = 6'h18 == s2_idx ? plru1_24 : _GEN_123; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_125 = 6'h19 == s2_idx ? plru1_25 : _GEN_124; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_126 = 6'h1a == s2_idx ? plru1_26 : _GEN_125; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_127 = 6'h1b == s2_idx ? plru1_27 : _GEN_126; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_128 = 6'h1c == s2_idx ? plru1_28 : _GEN_127; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_129 = 6'h1d == s2_idx ? plru1_29 : _GEN_128; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_130 = 6'h1e == s2_idx ? plru1_30 : _GEN_129; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_131 = 6'h1f == s2_idx ? plru1_31 : _GEN_130; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_132 = 6'h20 == s2_idx ? plru1_32 : _GEN_131; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_133 = 6'h21 == s2_idx ? plru1_33 : _GEN_132; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_134 = 6'h22 == s2_idx ? plru1_34 : _GEN_133; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_135 = 6'h23 == s2_idx ? plru1_35 : _GEN_134; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_136 = 6'h24 == s2_idx ? plru1_36 : _GEN_135; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_137 = 6'h25 == s2_idx ? plru1_37 : _GEN_136; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_138 = 6'h26 == s2_idx ? plru1_38 : _GEN_137; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_139 = 6'h27 == s2_idx ? plru1_39 : _GEN_138; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_140 = 6'h28 == s2_idx ? plru1_40 : _GEN_139; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_141 = 6'h29 == s2_idx ? plru1_41 : _GEN_140; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_142 = 6'h2a == s2_idx ? plru1_42 : _GEN_141; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_143 = 6'h2b == s2_idx ? plru1_43 : _GEN_142; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_144 = 6'h2c == s2_idx ? plru1_44 : _GEN_143; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_145 = 6'h2d == s2_idx ? plru1_45 : _GEN_144; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_146 = 6'h2e == s2_idx ? plru1_46 : _GEN_145; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_147 = 6'h2f == s2_idx ? plru1_47 : _GEN_146; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_148 = 6'h30 == s2_idx ? plru1_48 : _GEN_147; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_149 = 6'h31 == s2_idx ? plru1_49 : _GEN_148; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_150 = 6'h32 == s2_idx ? plru1_50 : _GEN_149; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_151 = 6'h33 == s2_idx ? plru1_51 : _GEN_150; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_152 = 6'h34 == s2_idx ? plru1_52 : _GEN_151; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_153 = 6'h35 == s2_idx ? plru1_53 : _GEN_152; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_154 = 6'h36 == s2_idx ? plru1_54 : _GEN_153; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_155 = 6'h37 == s2_idx ? plru1_55 : _GEN_154; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_156 = 6'h38 == s2_idx ? plru1_56 : _GEN_155; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_157 = 6'h39 == s2_idx ? plru1_57 : _GEN_156; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_158 = 6'h3a == s2_idx ? plru1_58 : _GEN_157; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_159 = 6'h3b == s2_idx ? plru1_59 : _GEN_158; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_160 = 6'h3c == s2_idx ? plru1_60 : _GEN_159; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_161 = 6'h3d == s2_idx ? plru1_61 : _GEN_160; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_162 = 6'h3e == s2_idx ? plru1_62 : _GEN_161; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_163 = 6'h3f == s2_idx ? plru1_63 : _GEN_162; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_165 = 6'h1 == s2_idx ? plru2_1 : plru2_0; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_166 = 6'h2 == s2_idx ? plru2_2 : _GEN_165; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_167 = 6'h3 == s2_idx ? plru2_3 : _GEN_166; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_168 = 6'h4 == s2_idx ? plru2_4 : _GEN_167; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_169 = 6'h5 == s2_idx ? plru2_5 : _GEN_168; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_170 = 6'h6 == s2_idx ? plru2_6 : _GEN_169; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_171 = 6'h7 == s2_idx ? plru2_7 : _GEN_170; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_172 = 6'h8 == s2_idx ? plru2_8 : _GEN_171; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_173 = 6'h9 == s2_idx ? plru2_9 : _GEN_172; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_174 = 6'ha == s2_idx ? plru2_10 : _GEN_173; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_175 = 6'hb == s2_idx ? plru2_11 : _GEN_174; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_176 = 6'hc == s2_idx ? plru2_12 : _GEN_175; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_177 = 6'hd == s2_idx ? plru2_13 : _GEN_176; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_178 = 6'he == s2_idx ? plru2_14 : _GEN_177; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_179 = 6'hf == s2_idx ? plru2_15 : _GEN_178; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_180 = 6'h10 == s2_idx ? plru2_16 : _GEN_179; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_181 = 6'h11 == s2_idx ? plru2_17 : _GEN_180; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_182 = 6'h12 == s2_idx ? plru2_18 : _GEN_181; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_183 = 6'h13 == s2_idx ? plru2_19 : _GEN_182; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_184 = 6'h14 == s2_idx ? plru2_20 : _GEN_183; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_185 = 6'h15 == s2_idx ? plru2_21 : _GEN_184; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_186 = 6'h16 == s2_idx ? plru2_22 : _GEN_185; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_187 = 6'h17 == s2_idx ? plru2_23 : _GEN_186; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_188 = 6'h18 == s2_idx ? plru2_24 : _GEN_187; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_189 = 6'h19 == s2_idx ? plru2_25 : _GEN_188; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_190 = 6'h1a == s2_idx ? plru2_26 : _GEN_189; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_191 = 6'h1b == s2_idx ? plru2_27 : _GEN_190; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_192 = 6'h1c == s2_idx ? plru2_28 : _GEN_191; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_193 = 6'h1d == s2_idx ? plru2_29 : _GEN_192; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_194 = 6'h1e == s2_idx ? plru2_30 : _GEN_193; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_195 = 6'h1f == s2_idx ? plru2_31 : _GEN_194; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_196 = 6'h20 == s2_idx ? plru2_32 : _GEN_195; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_197 = 6'h21 == s2_idx ? plru2_33 : _GEN_196; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_198 = 6'h22 == s2_idx ? plru2_34 : _GEN_197; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_199 = 6'h23 == s2_idx ? plru2_35 : _GEN_198; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_200 = 6'h24 == s2_idx ? plru2_36 : _GEN_199; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_201 = 6'h25 == s2_idx ? plru2_37 : _GEN_200; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_202 = 6'h26 == s2_idx ? plru2_38 : _GEN_201; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_203 = 6'h27 == s2_idx ? plru2_39 : _GEN_202; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_204 = 6'h28 == s2_idx ? plru2_40 : _GEN_203; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_205 = 6'h29 == s2_idx ? plru2_41 : _GEN_204; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_206 = 6'h2a == s2_idx ? plru2_42 : _GEN_205; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_207 = 6'h2b == s2_idx ? plru2_43 : _GEN_206; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_208 = 6'h2c == s2_idx ? plru2_44 : _GEN_207; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_209 = 6'h2d == s2_idx ? plru2_45 : _GEN_208; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_210 = 6'h2e == s2_idx ? plru2_46 : _GEN_209; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_211 = 6'h2f == s2_idx ? plru2_47 : _GEN_210; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_212 = 6'h30 == s2_idx ? plru2_48 : _GEN_211; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_213 = 6'h31 == s2_idx ? plru2_49 : _GEN_212; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_214 = 6'h32 == s2_idx ? plru2_50 : _GEN_213; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_215 = 6'h33 == s2_idx ? plru2_51 : _GEN_214; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_216 = 6'h34 == s2_idx ? plru2_52 : _GEN_215; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_217 = 6'h35 == s2_idx ? plru2_53 : _GEN_216; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_218 = 6'h36 == s2_idx ? plru2_54 : _GEN_217; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_219 = 6'h37 == s2_idx ? plru2_55 : _GEN_218; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_220 = 6'h38 == s2_idx ? plru2_56 : _GEN_219; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_221 = 6'h39 == s2_idx ? plru2_57 : _GEN_220; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_222 = 6'h3a == s2_idx ? plru2_58 : _GEN_221; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_223 = 6'h3b == s2_idx ? plru2_59 : _GEN_222; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_224 = 6'h3c == s2_idx ? plru2_60 : _GEN_223; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_225 = 6'h3d == s2_idx ? plru2_61 : _GEN_224; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_226 = 6'h3e == s2_idx ? plru2_62 : _GEN_225; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  _GEN_227 = 6'h3f == s2_idx ? plru2_63 : _GEN_226; // @[Cache.scala 256:25 Cache.scala 256:25]
  wire  replace_way_lo = ~_GEN_99 ? _GEN_163 : _GEN_227; // @[Cache.scala 256:25]
  wire [1:0] replace_way = {_GEN_99,replace_way_lo}; // @[Cat.scala 30:58]
  wire  dirty_out_0 = meta_0_io_dirty_r;
  wire  dirty_out_1 = meta_1_io_dirty_r;
  wire  _GEN_9 = 2'h1 == replace_way ? dirty_out_1 : dirty_out_0; // @[Cache.scala 250:18 Cache.scala 250:18]
  wire  dirty_out_2 = meta_2_io_dirty_r;
  wire  _GEN_10 = 2'h2 == replace_way ? dirty_out_2 : _GEN_9; // @[Cache.scala 250:18 Cache.scala 250:18]
  wire  dirty_out_3 = meta_3_io_dirty_r;
  wire [20:0] _GEN_13 = 2'h1 == replace_way ? tag_out_1 : tag_out_0; // @[Cache.scala 251:18 Cache.scala 251:18]
  wire [20:0] _GEN_14 = 2'h2 == replace_way ? tag_out_2 : _GEN_13; // @[Cache.scala 251:18 Cache.scala 251:18]
  wire [127:0] _GEN_17 = 2'h1 == replace_way ? sram_out_1 : sram_out_0; // @[Cache.scala 252:18 Cache.scala 252:18]
  wire [127:0] _GEN_18 = 2'h2 == replace_way ? sram_out_2 : _GEN_17; // @[Cache.scala 252:18 Cache.scala 252:18]
  wire  _GEN_27 = fi_ready ? io_in_req_bits_wen : s2_wen; // @[Cache.scala 238:24 Cache.scala 241:14 Cache.scala 213:25]
  reg [63:0] wdata1; // @[Cache.scala 258:23]
  reg [63:0] wdata2; // @[Cache.scala 259:23]
  wire  _T_2 = 4'h0 == state; // @[Conditional.scala 37:30]
  reg  REG_1; // @[Cache.scala 284:20]
  wire [63:0] _io_in_resp_bits_rdata_T_3 = s2_offs ? _GEN_7[127:64] : _GEN_7[63:0]; // @[Cache.scala 285:34]
  wire [63:0] _io_in_resp_bits_rdata_T_7 = s2_offs ? s2_reg_rdata[127:64] : s2_reg_rdata[63:0]; // @[Cache.scala 287:34]
  wire [63:0] _GEN_228 = REG_1 ? _io_in_resp_bits_rdata_T_3 : _io_in_resp_bits_rdata_T_7; // @[Cache.scala 284:37 Cache.scala 285:28 Cache.scala 287:28]
  reg  REG_2; // @[Cache.scala 289:20]
  wire  _plru0_T_1 = ~s2_way[1]; // @[Cache.scala 138:19]
  wire  _GEN_229 = 6'h0 == s2_idx ? ~s2_way[1] : plru0_0; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_230 = 6'h1 == s2_idx ? ~s2_way[1] : plru0_1; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_231 = 6'h2 == s2_idx ? ~s2_way[1] : plru0_2; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_232 = 6'h3 == s2_idx ? ~s2_way[1] : plru0_3; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_233 = 6'h4 == s2_idx ? ~s2_way[1] : plru0_4; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_234 = 6'h5 == s2_idx ? ~s2_way[1] : plru0_5; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_235 = 6'h6 == s2_idx ? ~s2_way[1] : plru0_6; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_236 = 6'h7 == s2_idx ? ~s2_way[1] : plru0_7; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_237 = 6'h8 == s2_idx ? ~s2_way[1] : plru0_8; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_238 = 6'h9 == s2_idx ? ~s2_way[1] : plru0_9; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_239 = 6'ha == s2_idx ? ~s2_way[1] : plru0_10; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_240 = 6'hb == s2_idx ? ~s2_way[1] : plru0_11; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_241 = 6'hc == s2_idx ? ~s2_way[1] : plru0_12; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_242 = 6'hd == s2_idx ? ~s2_way[1] : plru0_13; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_243 = 6'he == s2_idx ? ~s2_way[1] : plru0_14; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_244 = 6'hf == s2_idx ? ~s2_way[1] : plru0_15; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_245 = 6'h10 == s2_idx ? ~s2_way[1] : plru0_16; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_246 = 6'h11 == s2_idx ? ~s2_way[1] : plru0_17; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_247 = 6'h12 == s2_idx ? ~s2_way[1] : plru0_18; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_248 = 6'h13 == s2_idx ? ~s2_way[1] : plru0_19; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_249 = 6'h14 == s2_idx ? ~s2_way[1] : plru0_20; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_250 = 6'h15 == s2_idx ? ~s2_way[1] : plru0_21; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_251 = 6'h16 == s2_idx ? ~s2_way[1] : plru0_22; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_252 = 6'h17 == s2_idx ? ~s2_way[1] : plru0_23; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_253 = 6'h18 == s2_idx ? ~s2_way[1] : plru0_24; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_254 = 6'h19 == s2_idx ? ~s2_way[1] : plru0_25; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_255 = 6'h1a == s2_idx ? ~s2_way[1] : plru0_26; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_256 = 6'h1b == s2_idx ? ~s2_way[1] : plru0_27; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_257 = 6'h1c == s2_idx ? ~s2_way[1] : plru0_28; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_258 = 6'h1d == s2_idx ? ~s2_way[1] : plru0_29; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_259 = 6'h1e == s2_idx ? ~s2_way[1] : plru0_30; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_260 = 6'h1f == s2_idx ? ~s2_way[1] : plru0_31; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_261 = 6'h20 == s2_idx ? ~s2_way[1] : plru0_32; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_262 = 6'h21 == s2_idx ? ~s2_way[1] : plru0_33; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_263 = 6'h22 == s2_idx ? ~s2_way[1] : plru0_34; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_264 = 6'h23 == s2_idx ? ~s2_way[1] : plru0_35; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_265 = 6'h24 == s2_idx ? ~s2_way[1] : plru0_36; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_266 = 6'h25 == s2_idx ? ~s2_way[1] : plru0_37; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_267 = 6'h26 == s2_idx ? ~s2_way[1] : plru0_38; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_268 = 6'h27 == s2_idx ? ~s2_way[1] : plru0_39; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_269 = 6'h28 == s2_idx ? ~s2_way[1] : plru0_40; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_270 = 6'h29 == s2_idx ? ~s2_way[1] : plru0_41; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_271 = 6'h2a == s2_idx ? ~s2_way[1] : plru0_42; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_272 = 6'h2b == s2_idx ? ~s2_way[1] : plru0_43; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_273 = 6'h2c == s2_idx ? ~s2_way[1] : plru0_44; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_274 = 6'h2d == s2_idx ? ~s2_way[1] : plru0_45; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_275 = 6'h2e == s2_idx ? ~s2_way[1] : plru0_46; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_276 = 6'h2f == s2_idx ? ~s2_way[1] : plru0_47; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_277 = 6'h30 == s2_idx ? ~s2_way[1] : plru0_48; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_278 = 6'h31 == s2_idx ? ~s2_way[1] : plru0_49; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_279 = 6'h32 == s2_idx ? ~s2_way[1] : plru0_50; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_280 = 6'h33 == s2_idx ? ~s2_way[1] : plru0_51; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_281 = 6'h34 == s2_idx ? ~s2_way[1] : plru0_52; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_282 = 6'h35 == s2_idx ? ~s2_way[1] : plru0_53; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_283 = 6'h36 == s2_idx ? ~s2_way[1] : plru0_54; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_284 = 6'h37 == s2_idx ? ~s2_way[1] : plru0_55; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_285 = 6'h38 == s2_idx ? ~s2_way[1] : plru0_56; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_286 = 6'h39 == s2_idx ? ~s2_way[1] : plru0_57; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_287 = 6'h3a == s2_idx ? ~s2_way[1] : plru0_58; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_288 = 6'h3b == s2_idx ? ~s2_way[1] : plru0_59; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_289 = 6'h3c == s2_idx ? ~s2_way[1] : plru0_60; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_290 = 6'h3d == s2_idx ? ~s2_way[1] : plru0_61; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_291 = 6'h3e == s2_idx ? ~s2_way[1] : plru0_62; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_292 = 6'h3f == s2_idx ? ~s2_way[1] : plru0_63; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _plru1_T_1 = ~s2_way[0]; // @[Cache.scala 140:21]
  wire  _GEN_293 = 6'h0 == s2_idx ? ~s2_way[0] : plru1_0; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_294 = 6'h1 == s2_idx ? ~s2_way[0] : plru1_1; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_295 = 6'h2 == s2_idx ? ~s2_way[0] : plru1_2; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_296 = 6'h3 == s2_idx ? ~s2_way[0] : plru1_3; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_297 = 6'h4 == s2_idx ? ~s2_way[0] : plru1_4; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_298 = 6'h5 == s2_idx ? ~s2_way[0] : plru1_5; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_299 = 6'h6 == s2_idx ? ~s2_way[0] : plru1_6; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_300 = 6'h7 == s2_idx ? ~s2_way[0] : plru1_7; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_301 = 6'h8 == s2_idx ? ~s2_way[0] : plru1_8; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_302 = 6'h9 == s2_idx ? ~s2_way[0] : plru1_9; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_303 = 6'ha == s2_idx ? ~s2_way[0] : plru1_10; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_304 = 6'hb == s2_idx ? ~s2_way[0] : plru1_11; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_305 = 6'hc == s2_idx ? ~s2_way[0] : plru1_12; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_306 = 6'hd == s2_idx ? ~s2_way[0] : plru1_13; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_307 = 6'he == s2_idx ? ~s2_way[0] : plru1_14; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_308 = 6'hf == s2_idx ? ~s2_way[0] : plru1_15; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_309 = 6'h10 == s2_idx ? ~s2_way[0] : plru1_16; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_310 = 6'h11 == s2_idx ? ~s2_way[0] : plru1_17; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_311 = 6'h12 == s2_idx ? ~s2_way[0] : plru1_18; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_312 = 6'h13 == s2_idx ? ~s2_way[0] : plru1_19; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_313 = 6'h14 == s2_idx ? ~s2_way[0] : plru1_20; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_314 = 6'h15 == s2_idx ? ~s2_way[0] : plru1_21; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_315 = 6'h16 == s2_idx ? ~s2_way[0] : plru1_22; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_316 = 6'h17 == s2_idx ? ~s2_way[0] : plru1_23; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_317 = 6'h18 == s2_idx ? ~s2_way[0] : plru1_24; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_318 = 6'h19 == s2_idx ? ~s2_way[0] : plru1_25; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_319 = 6'h1a == s2_idx ? ~s2_way[0] : plru1_26; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_320 = 6'h1b == s2_idx ? ~s2_way[0] : plru1_27; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_321 = 6'h1c == s2_idx ? ~s2_way[0] : plru1_28; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_322 = 6'h1d == s2_idx ? ~s2_way[0] : plru1_29; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_323 = 6'h1e == s2_idx ? ~s2_way[0] : plru1_30; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_324 = 6'h1f == s2_idx ? ~s2_way[0] : plru1_31; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_325 = 6'h20 == s2_idx ? ~s2_way[0] : plru1_32; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_326 = 6'h21 == s2_idx ? ~s2_way[0] : plru1_33; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_327 = 6'h22 == s2_idx ? ~s2_way[0] : plru1_34; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_328 = 6'h23 == s2_idx ? ~s2_way[0] : plru1_35; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_329 = 6'h24 == s2_idx ? ~s2_way[0] : plru1_36; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_330 = 6'h25 == s2_idx ? ~s2_way[0] : plru1_37; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_331 = 6'h26 == s2_idx ? ~s2_way[0] : plru1_38; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_332 = 6'h27 == s2_idx ? ~s2_way[0] : plru1_39; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_333 = 6'h28 == s2_idx ? ~s2_way[0] : plru1_40; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_334 = 6'h29 == s2_idx ? ~s2_way[0] : plru1_41; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_335 = 6'h2a == s2_idx ? ~s2_way[0] : plru1_42; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_336 = 6'h2b == s2_idx ? ~s2_way[0] : plru1_43; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_337 = 6'h2c == s2_idx ? ~s2_way[0] : plru1_44; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_338 = 6'h2d == s2_idx ? ~s2_way[0] : plru1_45; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_339 = 6'h2e == s2_idx ? ~s2_way[0] : plru1_46; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_340 = 6'h2f == s2_idx ? ~s2_way[0] : plru1_47; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_341 = 6'h30 == s2_idx ? ~s2_way[0] : plru1_48; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_342 = 6'h31 == s2_idx ? ~s2_way[0] : plru1_49; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_343 = 6'h32 == s2_idx ? ~s2_way[0] : plru1_50; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_344 = 6'h33 == s2_idx ? ~s2_way[0] : plru1_51; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_345 = 6'h34 == s2_idx ? ~s2_way[0] : plru1_52; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_346 = 6'h35 == s2_idx ? ~s2_way[0] : plru1_53; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_347 = 6'h36 == s2_idx ? ~s2_way[0] : plru1_54; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_348 = 6'h37 == s2_idx ? ~s2_way[0] : plru1_55; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_349 = 6'h38 == s2_idx ? ~s2_way[0] : plru1_56; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_350 = 6'h39 == s2_idx ? ~s2_way[0] : plru1_57; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_351 = 6'h3a == s2_idx ? ~s2_way[0] : plru1_58; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_352 = 6'h3b == s2_idx ? ~s2_way[0] : plru1_59; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_353 = 6'h3c == s2_idx ? ~s2_way[0] : plru1_60; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_354 = 6'h3d == s2_idx ? ~s2_way[0] : plru1_61; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_355 = 6'h3e == s2_idx ? ~s2_way[0] : plru1_62; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_356 = 6'h3f == s2_idx ? ~s2_way[0] : plru1_63; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_357 = 6'h0 == s2_idx ? _plru1_T_1 : plru2_0; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_358 = 6'h1 == s2_idx ? _plru1_T_1 : plru2_1; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_359 = 6'h2 == s2_idx ? _plru1_T_1 : plru2_2; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_360 = 6'h3 == s2_idx ? _plru1_T_1 : plru2_3; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_361 = 6'h4 == s2_idx ? _plru1_T_1 : plru2_4; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_362 = 6'h5 == s2_idx ? _plru1_T_1 : plru2_5; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_363 = 6'h6 == s2_idx ? _plru1_T_1 : plru2_6; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_364 = 6'h7 == s2_idx ? _plru1_T_1 : plru2_7; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_365 = 6'h8 == s2_idx ? _plru1_T_1 : plru2_8; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_366 = 6'h9 == s2_idx ? _plru1_T_1 : plru2_9; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_367 = 6'ha == s2_idx ? _plru1_T_1 : plru2_10; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_368 = 6'hb == s2_idx ? _plru1_T_1 : plru2_11; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_369 = 6'hc == s2_idx ? _plru1_T_1 : plru2_12; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_370 = 6'hd == s2_idx ? _plru1_T_1 : plru2_13; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_371 = 6'he == s2_idx ? _plru1_T_1 : plru2_14; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_372 = 6'hf == s2_idx ? _plru1_T_1 : plru2_15; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_373 = 6'h10 == s2_idx ? _plru1_T_1 : plru2_16; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_374 = 6'h11 == s2_idx ? _plru1_T_1 : plru2_17; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_375 = 6'h12 == s2_idx ? _plru1_T_1 : plru2_18; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_376 = 6'h13 == s2_idx ? _plru1_T_1 : plru2_19; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_377 = 6'h14 == s2_idx ? _plru1_T_1 : plru2_20; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_378 = 6'h15 == s2_idx ? _plru1_T_1 : plru2_21; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_379 = 6'h16 == s2_idx ? _plru1_T_1 : plru2_22; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_380 = 6'h17 == s2_idx ? _plru1_T_1 : plru2_23; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_381 = 6'h18 == s2_idx ? _plru1_T_1 : plru2_24; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_382 = 6'h19 == s2_idx ? _plru1_T_1 : plru2_25; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_383 = 6'h1a == s2_idx ? _plru1_T_1 : plru2_26; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_384 = 6'h1b == s2_idx ? _plru1_T_1 : plru2_27; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_385 = 6'h1c == s2_idx ? _plru1_T_1 : plru2_28; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_386 = 6'h1d == s2_idx ? _plru1_T_1 : plru2_29; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_387 = 6'h1e == s2_idx ? _plru1_T_1 : plru2_30; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_388 = 6'h1f == s2_idx ? _plru1_T_1 : plru2_31; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_389 = 6'h20 == s2_idx ? _plru1_T_1 : plru2_32; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_390 = 6'h21 == s2_idx ? _plru1_T_1 : plru2_33; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_391 = 6'h22 == s2_idx ? _plru1_T_1 : plru2_34; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_392 = 6'h23 == s2_idx ? _plru1_T_1 : plru2_35; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_393 = 6'h24 == s2_idx ? _plru1_T_1 : plru2_36; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_394 = 6'h25 == s2_idx ? _plru1_T_1 : plru2_37; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_395 = 6'h26 == s2_idx ? _plru1_T_1 : plru2_38; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_396 = 6'h27 == s2_idx ? _plru1_T_1 : plru2_39; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_397 = 6'h28 == s2_idx ? _plru1_T_1 : plru2_40; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_398 = 6'h29 == s2_idx ? _plru1_T_1 : plru2_41; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_399 = 6'h2a == s2_idx ? _plru1_T_1 : plru2_42; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_400 = 6'h2b == s2_idx ? _plru1_T_1 : plru2_43; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_401 = 6'h2c == s2_idx ? _plru1_T_1 : plru2_44; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_402 = 6'h2d == s2_idx ? _plru1_T_1 : plru2_45; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_403 = 6'h2e == s2_idx ? _plru1_T_1 : plru2_46; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_404 = 6'h2f == s2_idx ? _plru1_T_1 : plru2_47; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_405 = 6'h30 == s2_idx ? _plru1_T_1 : plru2_48; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_406 = 6'h31 == s2_idx ? _plru1_T_1 : plru2_49; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_407 = 6'h32 == s2_idx ? _plru1_T_1 : plru2_50; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_408 = 6'h33 == s2_idx ? _plru1_T_1 : plru2_51; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_409 = 6'h34 == s2_idx ? _plru1_T_1 : plru2_52; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_410 = 6'h35 == s2_idx ? _plru1_T_1 : plru2_53; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_411 = 6'h36 == s2_idx ? _plru1_T_1 : plru2_54; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_412 = 6'h37 == s2_idx ? _plru1_T_1 : plru2_55; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_413 = 6'h38 == s2_idx ? _plru1_T_1 : plru2_56; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_414 = 6'h39 == s2_idx ? _plru1_T_1 : plru2_57; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_415 = 6'h3a == s2_idx ? _plru1_T_1 : plru2_58; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_416 = 6'h3b == s2_idx ? _plru1_T_1 : plru2_59; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_417 = 6'h3c == s2_idx ? _plru1_T_1 : plru2_60; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_418 = 6'h3d == s2_idx ? _plru1_T_1 : plru2_61; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_419 = 6'h3e == s2_idx ? _plru1_T_1 : plru2_62; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_420 = 6'h3f == s2_idx ? _plru1_T_1 : plru2_63; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_421 = _plru0_T_1 ? _GEN_293 : plru1_0; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_422 = _plru0_T_1 ? _GEN_294 : plru1_1; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_423 = _plru0_T_1 ? _GEN_295 : plru1_2; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_424 = _plru0_T_1 ? _GEN_296 : plru1_3; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_425 = _plru0_T_1 ? _GEN_297 : plru1_4; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_426 = _plru0_T_1 ? _GEN_298 : plru1_5; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_427 = _plru0_T_1 ? _GEN_299 : plru1_6; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_428 = _plru0_T_1 ? _GEN_300 : plru1_7; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_429 = _plru0_T_1 ? _GEN_301 : plru1_8; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_430 = _plru0_T_1 ? _GEN_302 : plru1_9; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_431 = _plru0_T_1 ? _GEN_303 : plru1_10; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_432 = _plru0_T_1 ? _GEN_304 : plru1_11; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_433 = _plru0_T_1 ? _GEN_305 : plru1_12; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_434 = _plru0_T_1 ? _GEN_306 : plru1_13; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_435 = _plru0_T_1 ? _GEN_307 : plru1_14; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_436 = _plru0_T_1 ? _GEN_308 : plru1_15; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_437 = _plru0_T_1 ? _GEN_309 : plru1_16; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_438 = _plru0_T_1 ? _GEN_310 : plru1_17; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_439 = _plru0_T_1 ? _GEN_311 : plru1_18; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_440 = _plru0_T_1 ? _GEN_312 : plru1_19; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_441 = _plru0_T_1 ? _GEN_313 : plru1_20; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_442 = _plru0_T_1 ? _GEN_314 : plru1_21; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_443 = _plru0_T_1 ? _GEN_315 : plru1_22; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_444 = _plru0_T_1 ? _GEN_316 : plru1_23; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_445 = _plru0_T_1 ? _GEN_317 : plru1_24; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_446 = _plru0_T_1 ? _GEN_318 : plru1_25; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_447 = _plru0_T_1 ? _GEN_319 : plru1_26; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_448 = _plru0_T_1 ? _GEN_320 : plru1_27; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_449 = _plru0_T_1 ? _GEN_321 : plru1_28; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_450 = _plru0_T_1 ? _GEN_322 : plru1_29; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_451 = _plru0_T_1 ? _GEN_323 : plru1_30; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_452 = _plru0_T_1 ? _GEN_324 : plru1_31; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_453 = _plru0_T_1 ? _GEN_325 : plru1_32; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_454 = _plru0_T_1 ? _GEN_326 : plru1_33; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_455 = _plru0_T_1 ? _GEN_327 : plru1_34; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_456 = _plru0_T_1 ? _GEN_328 : plru1_35; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_457 = _plru0_T_1 ? _GEN_329 : plru1_36; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_458 = _plru0_T_1 ? _GEN_330 : plru1_37; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_459 = _plru0_T_1 ? _GEN_331 : plru1_38; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_460 = _plru0_T_1 ? _GEN_332 : plru1_39; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_461 = _plru0_T_1 ? _GEN_333 : plru1_40; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_462 = _plru0_T_1 ? _GEN_334 : plru1_41; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_463 = _plru0_T_1 ? _GEN_335 : plru1_42; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_464 = _plru0_T_1 ? _GEN_336 : plru1_43; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_465 = _plru0_T_1 ? _GEN_337 : plru1_44; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_466 = _plru0_T_1 ? _GEN_338 : plru1_45; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_467 = _plru0_T_1 ? _GEN_339 : plru1_46; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_468 = _plru0_T_1 ? _GEN_340 : plru1_47; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_469 = _plru0_T_1 ? _GEN_341 : plru1_48; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_470 = _plru0_T_1 ? _GEN_342 : plru1_49; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_471 = _plru0_T_1 ? _GEN_343 : plru1_50; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_472 = _plru0_T_1 ? _GEN_344 : plru1_51; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_473 = _plru0_T_1 ? _GEN_345 : plru1_52; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_474 = _plru0_T_1 ? _GEN_346 : plru1_53; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_475 = _plru0_T_1 ? _GEN_347 : plru1_54; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_476 = _plru0_T_1 ? _GEN_348 : plru1_55; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_477 = _plru0_T_1 ? _GEN_349 : plru1_56; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_478 = _plru0_T_1 ? _GEN_350 : plru1_57; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_479 = _plru0_T_1 ? _GEN_351 : plru1_58; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_480 = _plru0_T_1 ? _GEN_352 : plru1_59; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_481 = _plru0_T_1 ? _GEN_353 : plru1_60; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_482 = _plru0_T_1 ? _GEN_354 : plru1_61; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_483 = _plru0_T_1 ? _GEN_355 : plru1_62; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_484 = _plru0_T_1 ? _GEN_356 : plru1_63; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_485 = _plru0_T_1 ? plru2_0 : _GEN_357; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_486 = _plru0_T_1 ? plru2_1 : _GEN_358; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_487 = _plru0_T_1 ? plru2_2 : _GEN_359; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_488 = _plru0_T_1 ? plru2_3 : _GEN_360; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_489 = _plru0_T_1 ? plru2_4 : _GEN_361; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_490 = _plru0_T_1 ? plru2_5 : _GEN_362; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_491 = _plru0_T_1 ? plru2_6 : _GEN_363; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_492 = _plru0_T_1 ? plru2_7 : _GEN_364; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_493 = _plru0_T_1 ? plru2_8 : _GEN_365; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_494 = _plru0_T_1 ? plru2_9 : _GEN_366; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_495 = _plru0_T_1 ? plru2_10 : _GEN_367; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_496 = _plru0_T_1 ? plru2_11 : _GEN_368; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_497 = _plru0_T_1 ? plru2_12 : _GEN_369; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_498 = _plru0_T_1 ? plru2_13 : _GEN_370; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_499 = _plru0_T_1 ? plru2_14 : _GEN_371; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_500 = _plru0_T_1 ? plru2_15 : _GEN_372; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_501 = _plru0_T_1 ? plru2_16 : _GEN_373; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_502 = _plru0_T_1 ? plru2_17 : _GEN_374; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_503 = _plru0_T_1 ? plru2_18 : _GEN_375; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_504 = _plru0_T_1 ? plru2_19 : _GEN_376; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_505 = _plru0_T_1 ? plru2_20 : _GEN_377; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_506 = _plru0_T_1 ? plru2_21 : _GEN_378; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_507 = _plru0_T_1 ? plru2_22 : _GEN_379; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_508 = _plru0_T_1 ? plru2_23 : _GEN_380; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_509 = _plru0_T_1 ? plru2_24 : _GEN_381; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_510 = _plru0_T_1 ? plru2_25 : _GEN_382; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_511 = _plru0_T_1 ? plru2_26 : _GEN_383; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_512 = _plru0_T_1 ? plru2_27 : _GEN_384; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_513 = _plru0_T_1 ? plru2_28 : _GEN_385; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_514 = _plru0_T_1 ? plru2_29 : _GEN_386; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_515 = _plru0_T_1 ? plru2_30 : _GEN_387; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_516 = _plru0_T_1 ? plru2_31 : _GEN_388; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_517 = _plru0_T_1 ? plru2_32 : _GEN_389; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_518 = _plru0_T_1 ? plru2_33 : _GEN_390; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_519 = _plru0_T_1 ? plru2_34 : _GEN_391; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_520 = _plru0_T_1 ? plru2_35 : _GEN_392; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_521 = _plru0_T_1 ? plru2_36 : _GEN_393; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_522 = _plru0_T_1 ? plru2_37 : _GEN_394; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_523 = _plru0_T_1 ? plru2_38 : _GEN_395; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_524 = _plru0_T_1 ? plru2_39 : _GEN_396; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_525 = _plru0_T_1 ? plru2_40 : _GEN_397; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_526 = _plru0_T_1 ? plru2_41 : _GEN_398; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_527 = _plru0_T_1 ? plru2_42 : _GEN_399; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_528 = _plru0_T_1 ? plru2_43 : _GEN_400; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_529 = _plru0_T_1 ? plru2_44 : _GEN_401; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_530 = _plru0_T_1 ? plru2_45 : _GEN_402; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_531 = _plru0_T_1 ? plru2_46 : _GEN_403; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_532 = _plru0_T_1 ? plru2_47 : _GEN_404; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_533 = _plru0_T_1 ? plru2_48 : _GEN_405; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_534 = _plru0_T_1 ? plru2_49 : _GEN_406; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_535 = _plru0_T_1 ? plru2_50 : _GEN_407; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_536 = _plru0_T_1 ? plru2_51 : _GEN_408; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_537 = _plru0_T_1 ? plru2_52 : _GEN_409; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_538 = _plru0_T_1 ? plru2_53 : _GEN_410; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_539 = _plru0_T_1 ? plru2_54 : _GEN_411; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_540 = _plru0_T_1 ? plru2_55 : _GEN_412; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_541 = _plru0_T_1 ? plru2_56 : _GEN_413; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_542 = _plru0_T_1 ? plru2_57 : _GEN_414; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_543 = _plru0_T_1 ? plru2_58 : _GEN_415; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_544 = _plru0_T_1 ? plru2_59 : _GEN_416; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_545 = _plru0_T_1 ? plru2_60 : _GEN_417; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_546 = _plru0_T_1 ? plru2_61 : _GEN_418; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_547 = _plru0_T_1 ? plru2_62 : _GEN_419; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_548 = _plru0_T_1 ? plru2_63 : _GEN_420; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _T_6 = s2_way == 2'h0; // @[Cache.scala 295:26]
  wire [7:0] sram_0_io_wdata_lo_lo_lo = s2_wmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] sram_0_io_wdata_lo_lo_hi = s2_wmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] sram_0_io_wdata_lo_hi_lo = s2_wmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] sram_0_io_wdata_lo_hi_hi = s2_wmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] sram_0_io_wdata_hi_lo_lo = s2_wmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] sram_0_io_wdata_hi_lo_hi = s2_wmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] sram_0_io_wdata_hi_hi_lo = s2_wmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] sram_0_io_wdata_hi_hi_hi = s2_wmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _sram_0_io_wdata_T_18 = {sram_0_io_wdata_hi_hi_hi,sram_0_io_wdata_hi_hi_lo,sram_0_io_wdata_hi_lo_hi,
    sram_0_io_wdata_hi_lo_lo,sram_0_io_wdata_lo_hi_hi,sram_0_io_wdata_lo_hi_lo,sram_0_io_wdata_lo_lo_hi,
    sram_0_io_wdata_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] _sram_0_io_wdata_T_19 = s2_wdata & _sram_0_io_wdata_T_18; // @[ID.scala 8:15]
  wire [63:0] _sram_0_io_wdata_T_20 = ~_sram_0_io_wdata_T_18; // @[ID.scala 8:37]
  wire [63:0] _sram_0_io_wdata_T_21 = _GEN_7[127:64] & _sram_0_io_wdata_T_20; // @[ID.scala 8:35]
  wire [63:0] sram_0_io_wdata_hi_1 = _sram_0_io_wdata_T_19 | _sram_0_io_wdata_T_21; // @[ID.scala 8:23]
  wire [127:0] _sram_0_io_wdata_T_22 = {sram_0_io_wdata_hi_1,_GEN_7[63:0]}; // @[Cat.scala 30:58]
  wire [63:0] _sram_0_io_wdata_T_43 = _GEN_7[63:0] & _sram_0_io_wdata_T_20; // @[ID.scala 8:35]
  wire [63:0] sram_0_io_wdata_lo_3 = _sram_0_io_wdata_T_19 | _sram_0_io_wdata_T_43; // @[ID.scala 8:23]
  wire [127:0] _sram_0_io_wdata_T_44 = {_GEN_7[127:64],sram_0_io_wdata_lo_3}; // @[Cat.scala 30:58]
  wire [127:0] _sram_0_io_wdata_T_45 = s2_offs ? _sram_0_io_wdata_T_22 : _sram_0_io_wdata_T_44; // @[Cache.scala 299:38]
  wire  _GEN_741 = s2_way == 2'h0 | fi_ready; // @[Cache.scala 295:35 Cache.scala 296:29]
  wire [5:0] _GEN_743 = s2_way == 2'h0 ? s2_idx : _GEN_3; // @[Cache.scala 295:35 Cache.scala 298:31]
  wire [127:0] _GEN_744 = s2_way == 2'h0 ? _sram_0_io_wdata_T_45 : 128'h0; // @[Cache.scala 295:35 Cache.scala 299:32 Cache.scala 112:16]
  wire  _T_7 = s2_way == 2'h1; // @[Cache.scala 295:26]
  wire  _GEN_745 = s2_way == 2'h1 | fi_ready; // @[Cache.scala 295:35 Cache.scala 296:29]
  wire [5:0] _GEN_747 = s2_way == 2'h1 ? s2_idx : _GEN_3; // @[Cache.scala 295:35 Cache.scala 298:31]
  wire [127:0] _GEN_748 = s2_way == 2'h1 ? _sram_0_io_wdata_T_45 : 128'h0; // @[Cache.scala 295:35 Cache.scala 299:32 Cache.scala 112:16]
  wire  _T_8 = s2_way == 2'h2; // @[Cache.scala 295:26]
  wire  _GEN_749 = s2_way == 2'h2 | fi_ready; // @[Cache.scala 295:35 Cache.scala 296:29]
  wire [5:0] _GEN_751 = s2_way == 2'h2 ? s2_idx : _GEN_3; // @[Cache.scala 295:35 Cache.scala 298:31]
  wire [127:0] _GEN_752 = s2_way == 2'h2 ? _sram_0_io_wdata_T_45 : 128'h0; // @[Cache.scala 295:35 Cache.scala 299:32 Cache.scala 112:16]
  wire  _T_9 = s2_way == 2'h3; // @[Cache.scala 295:26]
  wire  _GEN_753 = s2_way == 2'h3 | fi_ready; // @[Cache.scala 295:35 Cache.scala 296:29]
  wire [5:0] _GEN_755 = s2_way == 2'h3 ? s2_idx : _GEN_3; // @[Cache.scala 295:35 Cache.scala 298:31]
  wire [127:0] _GEN_756 = s2_way == 2'h3 ? _sram_0_io_wdata_T_45 : 128'h0; // @[Cache.scala 295:35 Cache.scala 299:32 Cache.scala 112:16]
  wire [3:0] _GEN_757 = ~s2_hit ? 4'h1 : state; // @[Cache.scala 308:31 Cache.scala 309:17 Cache.scala 207:22]
  wire  _GEN_758 = s2_hit & s2_wen ? _GEN_741 : fi_ready; // @[Cache.scala 293:33]
  wire  _GEN_759 = s2_hit & s2_wen & _T_6; // @[Cache.scala 293:33 Cache.scala 110:14]
  wire [5:0] _GEN_760 = s2_hit & s2_wen ? _GEN_743 : _GEN_3; // @[Cache.scala 293:33]
  wire [127:0] _GEN_761 = s2_hit & s2_wen ? _GEN_744 : 128'h0; // @[Cache.scala 293:33 Cache.scala 112:16]
  wire  _GEN_762 = s2_hit & s2_wen ? _GEN_745 : fi_ready; // @[Cache.scala 293:33]
  wire  _GEN_763 = s2_hit & s2_wen & _T_7; // @[Cache.scala 293:33 Cache.scala 110:14]
  wire [5:0] _GEN_764 = s2_hit & s2_wen ? _GEN_747 : _GEN_3; // @[Cache.scala 293:33]
  wire [127:0] _GEN_765 = s2_hit & s2_wen ? _GEN_748 : 128'h0; // @[Cache.scala 293:33 Cache.scala 112:16]
  wire  _GEN_766 = s2_hit & s2_wen ? _GEN_749 : fi_ready; // @[Cache.scala 293:33]
  wire  _GEN_767 = s2_hit & s2_wen & _T_8; // @[Cache.scala 293:33 Cache.scala 110:14]
  wire [5:0] _GEN_768 = s2_hit & s2_wen ? _GEN_751 : _GEN_3; // @[Cache.scala 293:33]
  wire [127:0] _GEN_769 = s2_hit & s2_wen ? _GEN_752 : 128'h0; // @[Cache.scala 293:33 Cache.scala 112:16]
  wire  _GEN_770 = s2_hit & s2_wen ? _GEN_753 : fi_ready; // @[Cache.scala 293:33]
  wire  _GEN_771 = s2_hit & s2_wen & _T_9; // @[Cache.scala 293:33 Cache.scala 110:14]
  wire [5:0] _GEN_772 = s2_hit & s2_wen ? _GEN_755 : _GEN_3; // @[Cache.scala 293:33]
  wire [127:0] _GEN_773 = s2_hit & s2_wen ? _GEN_756 : 128'h0; // @[Cache.scala 293:33 Cache.scala 112:16]
  wire [3:0] _GEN_774 = s2_hit & s2_wen ? 4'h7 : _GEN_757; // @[Cache.scala 293:33 Cache.scala 307:17]
  wire  _GEN_967 = REG_2 ? _GEN_758 : fi_ready; // @[Cache.scala 289:37]
  wire  _GEN_968 = REG_2 & _GEN_759; // @[Cache.scala 289:37 Cache.scala 110:14]
  wire [5:0] _GEN_969 = REG_2 ? _GEN_760 : _GEN_3; // @[Cache.scala 289:37]
  wire [127:0] _GEN_970 = REG_2 ? _GEN_761 : 128'h0; // @[Cache.scala 289:37 Cache.scala 112:16]
  wire  _GEN_971 = REG_2 ? _GEN_762 : fi_ready; // @[Cache.scala 289:37]
  wire  _GEN_972 = REG_2 & _GEN_763; // @[Cache.scala 289:37 Cache.scala 110:14]
  wire [5:0] _GEN_973 = REG_2 ? _GEN_764 : _GEN_3; // @[Cache.scala 289:37]
  wire [127:0] _GEN_974 = REG_2 ? _GEN_765 : 128'h0; // @[Cache.scala 289:37 Cache.scala 112:16]
  wire  _GEN_975 = REG_2 ? _GEN_766 : fi_ready; // @[Cache.scala 289:37]
  wire  _GEN_976 = REG_2 & _GEN_767; // @[Cache.scala 289:37 Cache.scala 110:14]
  wire [5:0] _GEN_977 = REG_2 ? _GEN_768 : _GEN_3; // @[Cache.scala 289:37]
  wire [127:0] _GEN_978 = REG_2 ? _GEN_769 : 128'h0; // @[Cache.scala 289:37 Cache.scala 112:16]
  wire  _GEN_979 = REG_2 ? _GEN_770 : fi_ready; // @[Cache.scala 289:37]
  wire  _GEN_980 = REG_2 & _GEN_771; // @[Cache.scala 289:37 Cache.scala 110:14]
  wire [5:0] _GEN_981 = REG_2 ? _GEN_772 : _GEN_3; // @[Cache.scala 289:37]
  wire [127:0] _GEN_982 = REG_2 ? _GEN_773 : 128'h0; // @[Cache.scala 289:37 Cache.scala 112:16]
  wire [3:0] _GEN_983 = REG_2 ? _GEN_774 : state; // @[Cache.scala 289:37 Cache.scala 207:22]
  wire  _T_11 = 4'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_984 = _T_12 ? 4'h2 : state; // @[Cache.scala 314:29 Cache.scala 315:15 Cache.scala 207:22]
  wire  _T_13 = 4'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_14 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_985 = ~io_out_resp_bits_rlast ? io_out_resp_bits_rdata : wdata1; // @[Cache.scala 320:37 Cache.scala 321:18 Cache.scala 258:23]
  wire [63:0] _GEN_986 = ~io_out_resp_bits_rlast ? wdata2 : io_out_resp_bits_rdata; // @[Cache.scala 320:37 Cache.scala 259:23 Cache.scala 323:18]
  wire [3:0] _GEN_987 = ~io_out_resp_bits_rlast ? state : 4'h3; // @[Cache.scala 320:37 Cache.scala 207:22 Cache.scala 324:17]
  wire [63:0] _GEN_988 = _T_14 ? _GEN_985 : wdata1; // @[Cache.scala 319:30 Cache.scala 258:23]
  wire [63:0] _GEN_989 = _T_14 ? _GEN_986 : wdata2; // @[Cache.scala 319:30 Cache.scala 259:23]
  wire [3:0] _GEN_990 = _T_14 ? _GEN_987 : state; // @[Cache.scala 319:30 Cache.scala 207:22]
  wire  _T_16 = 4'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_17 = replace_way == 2'h0; // @[Cache.scala 330:27]
  wire [63:0] _sram_0_io_wdata_T_66 = wdata2 & _sram_0_io_wdata_T_20; // @[ID.scala 8:35]
  wire [63:0] sram_0_io_wdata_hi_5 = _sram_0_io_wdata_T_19 | _sram_0_io_wdata_T_66; // @[ID.scala 8:23]
  wire [127:0] _sram_0_io_wdata_T_67 = {sram_0_io_wdata_hi_5,wdata1}; // @[Cat.scala 30:58]
  wire [63:0] _sram_0_io_wdata_T_87 = wdata1 & _sram_0_io_wdata_T_20; // @[ID.scala 8:35]
  wire [63:0] sram_0_io_wdata_lo_6 = _sram_0_io_wdata_T_19 | _sram_0_io_wdata_T_87; // @[ID.scala 8:23]
  wire [127:0] _sram_0_io_wdata_T_88 = {wdata2,sram_0_io_wdata_lo_6}; // @[Cat.scala 30:58]
  wire [127:0] _sram_0_io_wdata_T_89 = s2_offs ? _sram_0_io_wdata_T_67 : _sram_0_io_wdata_T_88; // @[Cache.scala 335:36]
  wire [127:0] _sram_0_io_wdata_T_90 = {wdata2,wdata1}; // @[Cat.scala 30:58]
  wire [127:0] _GEN_991 = s2_wen ? _sram_0_io_wdata_T_89 : _sram_0_io_wdata_T_90; // @[Cache.scala 334:25 Cache.scala 335:30 Cache.scala 339:30]
  wire  _GEN_992 = replace_way == 2'h0 | fi_ready; // @[Cache.scala 330:36 Cache.scala 331:25]
  wire [5:0] _GEN_994 = replace_way == 2'h0 ? s2_idx : _GEN_3; // @[Cache.scala 330:36 Cache.scala 333:27]
  wire [127:0] _GEN_995 = replace_way == 2'h0 ? _GEN_991 : 128'h0; // @[Cache.scala 330:36 Cache.scala 112:16]
  wire [20:0] _GEN_996 = replace_way == 2'h0 ? s2_tag : 21'h0; // @[Cache.scala 330:36 Cache.scala 344:28 Cache.scala 116:16]
  wire  _GEN_997 = replace_way == 2'h0 & s2_wen; // @[Cache.scala 330:36 Cache.scala 346:30 Cache.scala 118:18]
  wire  _T_18 = replace_way == 2'h1; // @[Cache.scala 330:27]
  wire  _GEN_999 = replace_way == 2'h1 | fi_ready; // @[Cache.scala 330:36 Cache.scala 331:25]
  wire [5:0] _GEN_1001 = replace_way == 2'h1 ? s2_idx : _GEN_3; // @[Cache.scala 330:36 Cache.scala 333:27]
  wire [127:0] _GEN_1002 = replace_way == 2'h1 ? _GEN_991 : 128'h0; // @[Cache.scala 330:36 Cache.scala 112:16]
  wire [20:0] _GEN_1003 = replace_way == 2'h1 ? s2_tag : 21'h0; // @[Cache.scala 330:36 Cache.scala 344:28 Cache.scala 116:16]
  wire  _GEN_1004 = replace_way == 2'h1 & s2_wen; // @[Cache.scala 330:36 Cache.scala 346:30 Cache.scala 118:18]
  wire  _T_19 = replace_way == 2'h2; // @[Cache.scala 330:27]
  wire  _GEN_1006 = replace_way == 2'h2 | fi_ready; // @[Cache.scala 330:36 Cache.scala 331:25]
  wire [5:0] _GEN_1008 = replace_way == 2'h2 ? s2_idx : _GEN_3; // @[Cache.scala 330:36 Cache.scala 333:27]
  wire [127:0] _GEN_1009 = replace_way == 2'h2 ? _GEN_991 : 128'h0; // @[Cache.scala 330:36 Cache.scala 112:16]
  wire [20:0] _GEN_1010 = replace_way == 2'h2 ? s2_tag : 21'h0; // @[Cache.scala 330:36 Cache.scala 344:28 Cache.scala 116:16]
  wire  _GEN_1011 = replace_way == 2'h2 & s2_wen; // @[Cache.scala 330:36 Cache.scala 346:30 Cache.scala 118:18]
  wire  _T_20 = replace_way == 2'h3; // @[Cache.scala 330:27]
  wire  _GEN_1013 = replace_way == 2'h3 | fi_ready; // @[Cache.scala 330:36 Cache.scala 331:25]
  wire [5:0] _GEN_1015 = replace_way == 2'h3 ? s2_idx : _GEN_3; // @[Cache.scala 330:36 Cache.scala 333:27]
  wire [127:0] _GEN_1016 = replace_way == 2'h3 ? _GEN_991 : 128'h0; // @[Cache.scala 330:36 Cache.scala 112:16]
  wire [20:0] _GEN_1017 = replace_way == 2'h3 ? s2_tag : 21'h0; // @[Cache.scala 330:36 Cache.scala 344:28 Cache.scala 116:16]
  wire  _GEN_1018 = replace_way == 2'h3 & s2_wen; // @[Cache.scala 330:36 Cache.scala 346:30 Cache.scala 118:18]
  wire  _plru0_T_3 = ~replace_way[1]; // @[Cache.scala 138:19]
  wire  _GEN_1019 = 6'h0 == s2_idx ? ~replace_way[1] : plru0_0; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1020 = 6'h1 == s2_idx ? ~replace_way[1] : plru0_1; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1021 = 6'h2 == s2_idx ? ~replace_way[1] : plru0_2; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1022 = 6'h3 == s2_idx ? ~replace_way[1] : plru0_3; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1023 = 6'h4 == s2_idx ? ~replace_way[1] : plru0_4; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1024 = 6'h5 == s2_idx ? ~replace_way[1] : plru0_5; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1025 = 6'h6 == s2_idx ? ~replace_way[1] : plru0_6; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1026 = 6'h7 == s2_idx ? ~replace_way[1] : plru0_7; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1027 = 6'h8 == s2_idx ? ~replace_way[1] : plru0_8; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1028 = 6'h9 == s2_idx ? ~replace_way[1] : plru0_9; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1029 = 6'ha == s2_idx ? ~replace_way[1] : plru0_10; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1030 = 6'hb == s2_idx ? ~replace_way[1] : plru0_11; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1031 = 6'hc == s2_idx ? ~replace_way[1] : plru0_12; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1032 = 6'hd == s2_idx ? ~replace_way[1] : plru0_13; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1033 = 6'he == s2_idx ? ~replace_way[1] : plru0_14; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1034 = 6'hf == s2_idx ? ~replace_way[1] : plru0_15; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1035 = 6'h10 == s2_idx ? ~replace_way[1] : plru0_16; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1036 = 6'h11 == s2_idx ? ~replace_way[1] : plru0_17; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1037 = 6'h12 == s2_idx ? ~replace_way[1] : plru0_18; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1038 = 6'h13 == s2_idx ? ~replace_way[1] : plru0_19; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1039 = 6'h14 == s2_idx ? ~replace_way[1] : plru0_20; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1040 = 6'h15 == s2_idx ? ~replace_way[1] : plru0_21; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1041 = 6'h16 == s2_idx ? ~replace_way[1] : plru0_22; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1042 = 6'h17 == s2_idx ? ~replace_way[1] : plru0_23; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1043 = 6'h18 == s2_idx ? ~replace_way[1] : plru0_24; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1044 = 6'h19 == s2_idx ? ~replace_way[1] : plru0_25; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1045 = 6'h1a == s2_idx ? ~replace_way[1] : plru0_26; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1046 = 6'h1b == s2_idx ? ~replace_way[1] : plru0_27; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1047 = 6'h1c == s2_idx ? ~replace_way[1] : plru0_28; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1048 = 6'h1d == s2_idx ? ~replace_way[1] : plru0_29; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1049 = 6'h1e == s2_idx ? ~replace_way[1] : plru0_30; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1050 = 6'h1f == s2_idx ? ~replace_way[1] : plru0_31; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1051 = 6'h20 == s2_idx ? ~replace_way[1] : plru0_32; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1052 = 6'h21 == s2_idx ? ~replace_way[1] : plru0_33; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1053 = 6'h22 == s2_idx ? ~replace_way[1] : plru0_34; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1054 = 6'h23 == s2_idx ? ~replace_way[1] : plru0_35; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1055 = 6'h24 == s2_idx ? ~replace_way[1] : plru0_36; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1056 = 6'h25 == s2_idx ? ~replace_way[1] : plru0_37; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1057 = 6'h26 == s2_idx ? ~replace_way[1] : plru0_38; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1058 = 6'h27 == s2_idx ? ~replace_way[1] : plru0_39; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1059 = 6'h28 == s2_idx ? ~replace_way[1] : plru0_40; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1060 = 6'h29 == s2_idx ? ~replace_way[1] : plru0_41; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1061 = 6'h2a == s2_idx ? ~replace_way[1] : plru0_42; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1062 = 6'h2b == s2_idx ? ~replace_way[1] : plru0_43; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1063 = 6'h2c == s2_idx ? ~replace_way[1] : plru0_44; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1064 = 6'h2d == s2_idx ? ~replace_way[1] : plru0_45; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1065 = 6'h2e == s2_idx ? ~replace_way[1] : plru0_46; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1066 = 6'h2f == s2_idx ? ~replace_way[1] : plru0_47; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1067 = 6'h30 == s2_idx ? ~replace_way[1] : plru0_48; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1068 = 6'h31 == s2_idx ? ~replace_way[1] : plru0_49; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1069 = 6'h32 == s2_idx ? ~replace_way[1] : plru0_50; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1070 = 6'h33 == s2_idx ? ~replace_way[1] : plru0_51; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1071 = 6'h34 == s2_idx ? ~replace_way[1] : plru0_52; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1072 = 6'h35 == s2_idx ? ~replace_way[1] : plru0_53; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1073 = 6'h36 == s2_idx ? ~replace_way[1] : plru0_54; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1074 = 6'h37 == s2_idx ? ~replace_way[1] : plru0_55; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1075 = 6'h38 == s2_idx ? ~replace_way[1] : plru0_56; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1076 = 6'h39 == s2_idx ? ~replace_way[1] : plru0_57; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1077 = 6'h3a == s2_idx ? ~replace_way[1] : plru0_58; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1078 = 6'h3b == s2_idx ? ~replace_way[1] : plru0_59; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1079 = 6'h3c == s2_idx ? ~replace_way[1] : plru0_60; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1080 = 6'h3d == s2_idx ? ~replace_way[1] : plru0_61; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1081 = 6'h3e == s2_idx ? ~replace_way[1] : plru0_62; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _GEN_1082 = 6'h3f == s2_idx ? ~replace_way[1] : plru0_63; // @[Cache.scala 138:16 Cache.scala 138:16 Cache.scala 131:22]
  wire  _plru1_T_3 = ~replace_way[0]; // @[Cache.scala 140:21]
  wire  _GEN_1083 = 6'h0 == s2_idx ? ~replace_way[0] : plru1_0; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1084 = 6'h1 == s2_idx ? ~replace_way[0] : plru1_1; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1085 = 6'h2 == s2_idx ? ~replace_way[0] : plru1_2; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1086 = 6'h3 == s2_idx ? ~replace_way[0] : plru1_3; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1087 = 6'h4 == s2_idx ? ~replace_way[0] : plru1_4; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1088 = 6'h5 == s2_idx ? ~replace_way[0] : plru1_5; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1089 = 6'h6 == s2_idx ? ~replace_way[0] : plru1_6; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1090 = 6'h7 == s2_idx ? ~replace_way[0] : plru1_7; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1091 = 6'h8 == s2_idx ? ~replace_way[0] : plru1_8; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1092 = 6'h9 == s2_idx ? ~replace_way[0] : plru1_9; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1093 = 6'ha == s2_idx ? ~replace_way[0] : plru1_10; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1094 = 6'hb == s2_idx ? ~replace_way[0] : plru1_11; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1095 = 6'hc == s2_idx ? ~replace_way[0] : plru1_12; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1096 = 6'hd == s2_idx ? ~replace_way[0] : plru1_13; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1097 = 6'he == s2_idx ? ~replace_way[0] : plru1_14; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1098 = 6'hf == s2_idx ? ~replace_way[0] : plru1_15; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1099 = 6'h10 == s2_idx ? ~replace_way[0] : plru1_16; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1100 = 6'h11 == s2_idx ? ~replace_way[0] : plru1_17; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1101 = 6'h12 == s2_idx ? ~replace_way[0] : plru1_18; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1102 = 6'h13 == s2_idx ? ~replace_way[0] : plru1_19; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1103 = 6'h14 == s2_idx ? ~replace_way[0] : plru1_20; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1104 = 6'h15 == s2_idx ? ~replace_way[0] : plru1_21; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1105 = 6'h16 == s2_idx ? ~replace_way[0] : plru1_22; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1106 = 6'h17 == s2_idx ? ~replace_way[0] : plru1_23; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1107 = 6'h18 == s2_idx ? ~replace_way[0] : plru1_24; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1108 = 6'h19 == s2_idx ? ~replace_way[0] : plru1_25; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1109 = 6'h1a == s2_idx ? ~replace_way[0] : plru1_26; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1110 = 6'h1b == s2_idx ? ~replace_way[0] : plru1_27; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1111 = 6'h1c == s2_idx ? ~replace_way[0] : plru1_28; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1112 = 6'h1d == s2_idx ? ~replace_way[0] : plru1_29; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1113 = 6'h1e == s2_idx ? ~replace_way[0] : plru1_30; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1114 = 6'h1f == s2_idx ? ~replace_way[0] : plru1_31; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1115 = 6'h20 == s2_idx ? ~replace_way[0] : plru1_32; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1116 = 6'h21 == s2_idx ? ~replace_way[0] : plru1_33; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1117 = 6'h22 == s2_idx ? ~replace_way[0] : plru1_34; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1118 = 6'h23 == s2_idx ? ~replace_way[0] : plru1_35; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1119 = 6'h24 == s2_idx ? ~replace_way[0] : plru1_36; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1120 = 6'h25 == s2_idx ? ~replace_way[0] : plru1_37; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1121 = 6'h26 == s2_idx ? ~replace_way[0] : plru1_38; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1122 = 6'h27 == s2_idx ? ~replace_way[0] : plru1_39; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1123 = 6'h28 == s2_idx ? ~replace_way[0] : plru1_40; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1124 = 6'h29 == s2_idx ? ~replace_way[0] : plru1_41; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1125 = 6'h2a == s2_idx ? ~replace_way[0] : plru1_42; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1126 = 6'h2b == s2_idx ? ~replace_way[0] : plru1_43; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1127 = 6'h2c == s2_idx ? ~replace_way[0] : plru1_44; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1128 = 6'h2d == s2_idx ? ~replace_way[0] : plru1_45; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1129 = 6'h2e == s2_idx ? ~replace_way[0] : plru1_46; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1130 = 6'h2f == s2_idx ? ~replace_way[0] : plru1_47; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1131 = 6'h30 == s2_idx ? ~replace_way[0] : plru1_48; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1132 = 6'h31 == s2_idx ? ~replace_way[0] : plru1_49; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1133 = 6'h32 == s2_idx ? ~replace_way[0] : plru1_50; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1134 = 6'h33 == s2_idx ? ~replace_way[0] : plru1_51; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1135 = 6'h34 == s2_idx ? ~replace_way[0] : plru1_52; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1136 = 6'h35 == s2_idx ? ~replace_way[0] : plru1_53; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1137 = 6'h36 == s2_idx ? ~replace_way[0] : plru1_54; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1138 = 6'h37 == s2_idx ? ~replace_way[0] : plru1_55; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1139 = 6'h38 == s2_idx ? ~replace_way[0] : plru1_56; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1140 = 6'h39 == s2_idx ? ~replace_way[0] : plru1_57; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1141 = 6'h3a == s2_idx ? ~replace_way[0] : plru1_58; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1142 = 6'h3b == s2_idx ? ~replace_way[0] : plru1_59; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1143 = 6'h3c == s2_idx ? ~replace_way[0] : plru1_60; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1144 = 6'h3d == s2_idx ? ~replace_way[0] : plru1_61; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1145 = 6'h3e == s2_idx ? ~replace_way[0] : plru1_62; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1146 = 6'h3f == s2_idx ? ~replace_way[0] : plru1_63; // @[Cache.scala 140:18 Cache.scala 140:18 Cache.scala 133:22]
  wire  _GEN_1147 = 6'h0 == s2_idx ? _plru1_T_3 : plru2_0; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1148 = 6'h1 == s2_idx ? _plru1_T_3 : plru2_1; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1149 = 6'h2 == s2_idx ? _plru1_T_3 : plru2_2; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1150 = 6'h3 == s2_idx ? _plru1_T_3 : plru2_3; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1151 = 6'h4 == s2_idx ? _plru1_T_3 : plru2_4; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1152 = 6'h5 == s2_idx ? _plru1_T_3 : plru2_5; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1153 = 6'h6 == s2_idx ? _plru1_T_3 : plru2_6; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1154 = 6'h7 == s2_idx ? _plru1_T_3 : plru2_7; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1155 = 6'h8 == s2_idx ? _plru1_T_3 : plru2_8; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1156 = 6'h9 == s2_idx ? _plru1_T_3 : plru2_9; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1157 = 6'ha == s2_idx ? _plru1_T_3 : plru2_10; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1158 = 6'hb == s2_idx ? _plru1_T_3 : plru2_11; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1159 = 6'hc == s2_idx ? _plru1_T_3 : plru2_12; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1160 = 6'hd == s2_idx ? _plru1_T_3 : plru2_13; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1161 = 6'he == s2_idx ? _plru1_T_3 : plru2_14; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1162 = 6'hf == s2_idx ? _plru1_T_3 : plru2_15; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1163 = 6'h10 == s2_idx ? _plru1_T_3 : plru2_16; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1164 = 6'h11 == s2_idx ? _plru1_T_3 : plru2_17; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1165 = 6'h12 == s2_idx ? _plru1_T_3 : plru2_18; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1166 = 6'h13 == s2_idx ? _plru1_T_3 : plru2_19; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1167 = 6'h14 == s2_idx ? _plru1_T_3 : plru2_20; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1168 = 6'h15 == s2_idx ? _plru1_T_3 : plru2_21; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1169 = 6'h16 == s2_idx ? _plru1_T_3 : plru2_22; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1170 = 6'h17 == s2_idx ? _plru1_T_3 : plru2_23; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1171 = 6'h18 == s2_idx ? _plru1_T_3 : plru2_24; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1172 = 6'h19 == s2_idx ? _plru1_T_3 : plru2_25; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1173 = 6'h1a == s2_idx ? _plru1_T_3 : plru2_26; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1174 = 6'h1b == s2_idx ? _plru1_T_3 : plru2_27; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1175 = 6'h1c == s2_idx ? _plru1_T_3 : plru2_28; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1176 = 6'h1d == s2_idx ? _plru1_T_3 : plru2_29; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1177 = 6'h1e == s2_idx ? _plru1_T_3 : plru2_30; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1178 = 6'h1f == s2_idx ? _plru1_T_3 : plru2_31; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1179 = 6'h20 == s2_idx ? _plru1_T_3 : plru2_32; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1180 = 6'h21 == s2_idx ? _plru1_T_3 : plru2_33; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1181 = 6'h22 == s2_idx ? _plru1_T_3 : plru2_34; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1182 = 6'h23 == s2_idx ? _plru1_T_3 : plru2_35; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1183 = 6'h24 == s2_idx ? _plru1_T_3 : plru2_36; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1184 = 6'h25 == s2_idx ? _plru1_T_3 : plru2_37; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1185 = 6'h26 == s2_idx ? _plru1_T_3 : plru2_38; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1186 = 6'h27 == s2_idx ? _plru1_T_3 : plru2_39; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1187 = 6'h28 == s2_idx ? _plru1_T_3 : plru2_40; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1188 = 6'h29 == s2_idx ? _plru1_T_3 : plru2_41; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1189 = 6'h2a == s2_idx ? _plru1_T_3 : plru2_42; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1190 = 6'h2b == s2_idx ? _plru1_T_3 : plru2_43; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1191 = 6'h2c == s2_idx ? _plru1_T_3 : plru2_44; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1192 = 6'h2d == s2_idx ? _plru1_T_3 : plru2_45; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1193 = 6'h2e == s2_idx ? _plru1_T_3 : plru2_46; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1194 = 6'h2f == s2_idx ? _plru1_T_3 : plru2_47; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1195 = 6'h30 == s2_idx ? _plru1_T_3 : plru2_48; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1196 = 6'h31 == s2_idx ? _plru1_T_3 : plru2_49; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1197 = 6'h32 == s2_idx ? _plru1_T_3 : plru2_50; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1198 = 6'h33 == s2_idx ? _plru1_T_3 : plru2_51; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1199 = 6'h34 == s2_idx ? _plru1_T_3 : plru2_52; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1200 = 6'h35 == s2_idx ? _plru1_T_3 : plru2_53; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1201 = 6'h36 == s2_idx ? _plru1_T_3 : plru2_54; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1202 = 6'h37 == s2_idx ? _plru1_T_3 : plru2_55; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1203 = 6'h38 == s2_idx ? _plru1_T_3 : plru2_56; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1204 = 6'h39 == s2_idx ? _plru1_T_3 : plru2_57; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1205 = 6'h3a == s2_idx ? _plru1_T_3 : plru2_58; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1206 = 6'h3b == s2_idx ? _plru1_T_3 : plru2_59; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1207 = 6'h3c == s2_idx ? _plru1_T_3 : plru2_60; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1208 = 6'h3d == s2_idx ? _plru1_T_3 : plru2_61; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1209 = 6'h3e == s2_idx ? _plru1_T_3 : plru2_62; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1210 = 6'h3f == s2_idx ? _plru1_T_3 : plru2_63; // @[Cache.scala 142:18 Cache.scala 142:18 Cache.scala 135:22]
  wire  _GEN_1211 = _plru0_T_3 ? _GEN_1083 : plru1_0; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1212 = _plru0_T_3 ? _GEN_1084 : plru1_1; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1213 = _plru0_T_3 ? _GEN_1085 : plru1_2; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1214 = _plru0_T_3 ? _GEN_1086 : plru1_3; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1215 = _plru0_T_3 ? _GEN_1087 : plru1_4; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1216 = _plru0_T_3 ? _GEN_1088 : plru1_5; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1217 = _plru0_T_3 ? _GEN_1089 : plru1_6; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1218 = _plru0_T_3 ? _GEN_1090 : plru1_7; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1219 = _plru0_T_3 ? _GEN_1091 : plru1_8; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1220 = _plru0_T_3 ? _GEN_1092 : plru1_9; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1221 = _plru0_T_3 ? _GEN_1093 : plru1_10; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1222 = _plru0_T_3 ? _GEN_1094 : plru1_11; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1223 = _plru0_T_3 ? _GEN_1095 : plru1_12; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1224 = _plru0_T_3 ? _GEN_1096 : plru1_13; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1225 = _plru0_T_3 ? _GEN_1097 : plru1_14; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1226 = _plru0_T_3 ? _GEN_1098 : plru1_15; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1227 = _plru0_T_3 ? _GEN_1099 : plru1_16; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1228 = _plru0_T_3 ? _GEN_1100 : plru1_17; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1229 = _plru0_T_3 ? _GEN_1101 : plru1_18; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1230 = _plru0_T_3 ? _GEN_1102 : plru1_19; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1231 = _plru0_T_3 ? _GEN_1103 : plru1_20; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1232 = _plru0_T_3 ? _GEN_1104 : plru1_21; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1233 = _plru0_T_3 ? _GEN_1105 : plru1_22; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1234 = _plru0_T_3 ? _GEN_1106 : plru1_23; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1235 = _plru0_T_3 ? _GEN_1107 : plru1_24; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1236 = _plru0_T_3 ? _GEN_1108 : plru1_25; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1237 = _plru0_T_3 ? _GEN_1109 : plru1_26; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1238 = _plru0_T_3 ? _GEN_1110 : plru1_27; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1239 = _plru0_T_3 ? _GEN_1111 : plru1_28; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1240 = _plru0_T_3 ? _GEN_1112 : plru1_29; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1241 = _plru0_T_3 ? _GEN_1113 : plru1_30; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1242 = _plru0_T_3 ? _GEN_1114 : plru1_31; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1243 = _plru0_T_3 ? _GEN_1115 : plru1_32; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1244 = _plru0_T_3 ? _GEN_1116 : plru1_33; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1245 = _plru0_T_3 ? _GEN_1117 : plru1_34; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1246 = _plru0_T_3 ? _GEN_1118 : plru1_35; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1247 = _plru0_T_3 ? _GEN_1119 : plru1_36; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1248 = _plru0_T_3 ? _GEN_1120 : plru1_37; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1249 = _plru0_T_3 ? _GEN_1121 : plru1_38; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1250 = _plru0_T_3 ? _GEN_1122 : plru1_39; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1251 = _plru0_T_3 ? _GEN_1123 : plru1_40; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1252 = _plru0_T_3 ? _GEN_1124 : plru1_41; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1253 = _plru0_T_3 ? _GEN_1125 : plru1_42; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1254 = _plru0_T_3 ? _GEN_1126 : plru1_43; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1255 = _plru0_T_3 ? _GEN_1127 : plru1_44; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1256 = _plru0_T_3 ? _GEN_1128 : plru1_45; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1257 = _plru0_T_3 ? _GEN_1129 : plru1_46; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1258 = _plru0_T_3 ? _GEN_1130 : plru1_47; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1259 = _plru0_T_3 ? _GEN_1131 : plru1_48; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1260 = _plru0_T_3 ? _GEN_1132 : plru1_49; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1261 = _plru0_T_3 ? _GEN_1133 : plru1_50; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1262 = _plru0_T_3 ? _GEN_1134 : plru1_51; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1263 = _plru0_T_3 ? _GEN_1135 : plru1_52; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1264 = _plru0_T_3 ? _GEN_1136 : plru1_53; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1265 = _plru0_T_3 ? _GEN_1137 : plru1_54; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1266 = _plru0_T_3 ? _GEN_1138 : plru1_55; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1267 = _plru0_T_3 ? _GEN_1139 : plru1_56; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1268 = _plru0_T_3 ? _GEN_1140 : plru1_57; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1269 = _plru0_T_3 ? _GEN_1141 : plru1_58; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1270 = _plru0_T_3 ? _GEN_1142 : plru1_59; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1271 = _plru0_T_3 ? _GEN_1143 : plru1_60; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1272 = _plru0_T_3 ? _GEN_1144 : plru1_61; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1273 = _plru0_T_3 ? _GEN_1145 : plru1_62; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1274 = _plru0_T_3 ? _GEN_1146 : plru1_63; // @[Cache.scala 139:27 Cache.scala 133:22]
  wire  _GEN_1275 = _plru0_T_3 ? plru2_0 : _GEN_1147; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1276 = _plru0_T_3 ? plru2_1 : _GEN_1148; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1277 = _plru0_T_3 ? plru2_2 : _GEN_1149; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1278 = _plru0_T_3 ? plru2_3 : _GEN_1150; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1279 = _plru0_T_3 ? plru2_4 : _GEN_1151; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1280 = _plru0_T_3 ? plru2_5 : _GEN_1152; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1281 = _plru0_T_3 ? plru2_6 : _GEN_1153; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1282 = _plru0_T_3 ? plru2_7 : _GEN_1154; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1283 = _plru0_T_3 ? plru2_8 : _GEN_1155; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1284 = _plru0_T_3 ? plru2_9 : _GEN_1156; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1285 = _plru0_T_3 ? plru2_10 : _GEN_1157; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1286 = _plru0_T_3 ? plru2_11 : _GEN_1158; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1287 = _plru0_T_3 ? plru2_12 : _GEN_1159; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1288 = _plru0_T_3 ? plru2_13 : _GEN_1160; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1289 = _plru0_T_3 ? plru2_14 : _GEN_1161; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1290 = _plru0_T_3 ? plru2_15 : _GEN_1162; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1291 = _plru0_T_3 ? plru2_16 : _GEN_1163; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1292 = _plru0_T_3 ? plru2_17 : _GEN_1164; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1293 = _plru0_T_3 ? plru2_18 : _GEN_1165; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1294 = _plru0_T_3 ? plru2_19 : _GEN_1166; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1295 = _plru0_T_3 ? plru2_20 : _GEN_1167; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1296 = _plru0_T_3 ? plru2_21 : _GEN_1168; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1297 = _plru0_T_3 ? plru2_22 : _GEN_1169; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1298 = _plru0_T_3 ? plru2_23 : _GEN_1170; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1299 = _plru0_T_3 ? plru2_24 : _GEN_1171; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1300 = _plru0_T_3 ? plru2_25 : _GEN_1172; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1301 = _plru0_T_3 ? plru2_26 : _GEN_1173; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1302 = _plru0_T_3 ? plru2_27 : _GEN_1174; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1303 = _plru0_T_3 ? plru2_28 : _GEN_1175; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1304 = _plru0_T_3 ? plru2_29 : _GEN_1176; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1305 = _plru0_T_3 ? plru2_30 : _GEN_1177; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1306 = _plru0_T_3 ? plru2_31 : _GEN_1178; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1307 = _plru0_T_3 ? plru2_32 : _GEN_1179; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1308 = _plru0_T_3 ? plru2_33 : _GEN_1180; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1309 = _plru0_T_3 ? plru2_34 : _GEN_1181; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1310 = _plru0_T_3 ? plru2_35 : _GEN_1182; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1311 = _plru0_T_3 ? plru2_36 : _GEN_1183; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1312 = _plru0_T_3 ? plru2_37 : _GEN_1184; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1313 = _plru0_T_3 ? plru2_38 : _GEN_1185; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1314 = _plru0_T_3 ? plru2_39 : _GEN_1186; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1315 = _plru0_T_3 ? plru2_40 : _GEN_1187; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1316 = _plru0_T_3 ? plru2_41 : _GEN_1188; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1317 = _plru0_T_3 ? plru2_42 : _GEN_1189; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1318 = _plru0_T_3 ? plru2_43 : _GEN_1190; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1319 = _plru0_T_3 ? plru2_44 : _GEN_1191; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1320 = _plru0_T_3 ? plru2_45 : _GEN_1192; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1321 = _plru0_T_3 ? plru2_46 : _GEN_1193; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1322 = _plru0_T_3 ? plru2_47 : _GEN_1194; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1323 = _plru0_T_3 ? plru2_48 : _GEN_1195; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1324 = _plru0_T_3 ? plru2_49 : _GEN_1196; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1325 = _plru0_T_3 ? plru2_50 : _GEN_1197; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1326 = _plru0_T_3 ? plru2_51 : _GEN_1198; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1327 = _plru0_T_3 ? plru2_52 : _GEN_1199; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1328 = _plru0_T_3 ? plru2_53 : _GEN_1200; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1329 = _plru0_T_3 ? plru2_54 : _GEN_1201; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1330 = _plru0_T_3 ? plru2_55 : _GEN_1202; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1331 = _plru0_T_3 ? plru2_56 : _GEN_1203; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1332 = _plru0_T_3 ? plru2_57 : _GEN_1204; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1333 = _plru0_T_3 ? plru2_58 : _GEN_1205; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1334 = _plru0_T_3 ? plru2_59 : _GEN_1206; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1335 = _plru0_T_3 ? plru2_60 : _GEN_1207; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1336 = _plru0_T_3 ? plru2_61 : _GEN_1208; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1337 = _plru0_T_3 ? plru2_62 : _GEN_1209; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire  _GEN_1338 = _plru0_T_3 ? plru2_63 : _GEN_1210; // @[Cache.scala 139:27 Cache.scala 135:22]
  wire [3:0] _GEN_1339 = s2_reg_dirty ? 4'h4 : 4'h7; // @[Cache.scala 349:27 Cache.scala 350:15 Cache.scala 353:15]
  wire  _GEN_1340 = s2_reg_dirty ? plru0_0 : _GEN_1019; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1341 = s2_reg_dirty ? plru0_1 : _GEN_1020; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1342 = s2_reg_dirty ? plru0_2 : _GEN_1021; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1343 = s2_reg_dirty ? plru0_3 : _GEN_1022; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1344 = s2_reg_dirty ? plru0_4 : _GEN_1023; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1345 = s2_reg_dirty ? plru0_5 : _GEN_1024; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1346 = s2_reg_dirty ? plru0_6 : _GEN_1025; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1347 = s2_reg_dirty ? plru0_7 : _GEN_1026; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1348 = s2_reg_dirty ? plru0_8 : _GEN_1027; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1349 = s2_reg_dirty ? plru0_9 : _GEN_1028; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1350 = s2_reg_dirty ? plru0_10 : _GEN_1029; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1351 = s2_reg_dirty ? plru0_11 : _GEN_1030; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1352 = s2_reg_dirty ? plru0_12 : _GEN_1031; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1353 = s2_reg_dirty ? plru0_13 : _GEN_1032; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1354 = s2_reg_dirty ? plru0_14 : _GEN_1033; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1355 = s2_reg_dirty ? plru0_15 : _GEN_1034; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1356 = s2_reg_dirty ? plru0_16 : _GEN_1035; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1357 = s2_reg_dirty ? plru0_17 : _GEN_1036; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1358 = s2_reg_dirty ? plru0_18 : _GEN_1037; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1359 = s2_reg_dirty ? plru0_19 : _GEN_1038; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1360 = s2_reg_dirty ? plru0_20 : _GEN_1039; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1361 = s2_reg_dirty ? plru0_21 : _GEN_1040; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1362 = s2_reg_dirty ? plru0_22 : _GEN_1041; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1363 = s2_reg_dirty ? plru0_23 : _GEN_1042; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1364 = s2_reg_dirty ? plru0_24 : _GEN_1043; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1365 = s2_reg_dirty ? plru0_25 : _GEN_1044; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1366 = s2_reg_dirty ? plru0_26 : _GEN_1045; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1367 = s2_reg_dirty ? plru0_27 : _GEN_1046; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1368 = s2_reg_dirty ? plru0_28 : _GEN_1047; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1369 = s2_reg_dirty ? plru0_29 : _GEN_1048; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1370 = s2_reg_dirty ? plru0_30 : _GEN_1049; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1371 = s2_reg_dirty ? plru0_31 : _GEN_1050; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1372 = s2_reg_dirty ? plru0_32 : _GEN_1051; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1373 = s2_reg_dirty ? plru0_33 : _GEN_1052; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1374 = s2_reg_dirty ? plru0_34 : _GEN_1053; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1375 = s2_reg_dirty ? plru0_35 : _GEN_1054; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1376 = s2_reg_dirty ? plru0_36 : _GEN_1055; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1377 = s2_reg_dirty ? plru0_37 : _GEN_1056; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1378 = s2_reg_dirty ? plru0_38 : _GEN_1057; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1379 = s2_reg_dirty ? plru0_39 : _GEN_1058; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1380 = s2_reg_dirty ? plru0_40 : _GEN_1059; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1381 = s2_reg_dirty ? plru0_41 : _GEN_1060; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1382 = s2_reg_dirty ? plru0_42 : _GEN_1061; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1383 = s2_reg_dirty ? plru0_43 : _GEN_1062; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1384 = s2_reg_dirty ? plru0_44 : _GEN_1063; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1385 = s2_reg_dirty ? plru0_45 : _GEN_1064; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1386 = s2_reg_dirty ? plru0_46 : _GEN_1065; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1387 = s2_reg_dirty ? plru0_47 : _GEN_1066; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1388 = s2_reg_dirty ? plru0_48 : _GEN_1067; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1389 = s2_reg_dirty ? plru0_49 : _GEN_1068; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1390 = s2_reg_dirty ? plru0_50 : _GEN_1069; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1391 = s2_reg_dirty ? plru0_51 : _GEN_1070; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1392 = s2_reg_dirty ? plru0_52 : _GEN_1071; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1393 = s2_reg_dirty ? plru0_53 : _GEN_1072; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1394 = s2_reg_dirty ? plru0_54 : _GEN_1073; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1395 = s2_reg_dirty ? plru0_55 : _GEN_1074; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1396 = s2_reg_dirty ? plru0_56 : _GEN_1075; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1397 = s2_reg_dirty ? plru0_57 : _GEN_1076; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1398 = s2_reg_dirty ? plru0_58 : _GEN_1077; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1399 = s2_reg_dirty ? plru0_59 : _GEN_1078; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1400 = s2_reg_dirty ? plru0_60 : _GEN_1079; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1401 = s2_reg_dirty ? plru0_61 : _GEN_1080; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1402 = s2_reg_dirty ? plru0_62 : _GEN_1081; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1403 = s2_reg_dirty ? plru0_63 : _GEN_1082; // @[Cache.scala 349:27 Cache.scala 131:22]
  wire  _GEN_1404 = s2_reg_dirty ? plru1_0 : _GEN_1211; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1405 = s2_reg_dirty ? plru1_1 : _GEN_1212; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1406 = s2_reg_dirty ? plru1_2 : _GEN_1213; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1407 = s2_reg_dirty ? plru1_3 : _GEN_1214; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1408 = s2_reg_dirty ? plru1_4 : _GEN_1215; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1409 = s2_reg_dirty ? plru1_5 : _GEN_1216; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1410 = s2_reg_dirty ? plru1_6 : _GEN_1217; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1411 = s2_reg_dirty ? plru1_7 : _GEN_1218; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1412 = s2_reg_dirty ? plru1_8 : _GEN_1219; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1413 = s2_reg_dirty ? plru1_9 : _GEN_1220; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1414 = s2_reg_dirty ? plru1_10 : _GEN_1221; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1415 = s2_reg_dirty ? plru1_11 : _GEN_1222; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1416 = s2_reg_dirty ? plru1_12 : _GEN_1223; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1417 = s2_reg_dirty ? plru1_13 : _GEN_1224; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1418 = s2_reg_dirty ? plru1_14 : _GEN_1225; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1419 = s2_reg_dirty ? plru1_15 : _GEN_1226; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1420 = s2_reg_dirty ? plru1_16 : _GEN_1227; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1421 = s2_reg_dirty ? plru1_17 : _GEN_1228; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1422 = s2_reg_dirty ? plru1_18 : _GEN_1229; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1423 = s2_reg_dirty ? plru1_19 : _GEN_1230; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1424 = s2_reg_dirty ? plru1_20 : _GEN_1231; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1425 = s2_reg_dirty ? plru1_21 : _GEN_1232; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1426 = s2_reg_dirty ? plru1_22 : _GEN_1233; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1427 = s2_reg_dirty ? plru1_23 : _GEN_1234; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1428 = s2_reg_dirty ? plru1_24 : _GEN_1235; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1429 = s2_reg_dirty ? plru1_25 : _GEN_1236; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1430 = s2_reg_dirty ? plru1_26 : _GEN_1237; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1431 = s2_reg_dirty ? plru1_27 : _GEN_1238; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1432 = s2_reg_dirty ? plru1_28 : _GEN_1239; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1433 = s2_reg_dirty ? plru1_29 : _GEN_1240; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1434 = s2_reg_dirty ? plru1_30 : _GEN_1241; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1435 = s2_reg_dirty ? plru1_31 : _GEN_1242; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1436 = s2_reg_dirty ? plru1_32 : _GEN_1243; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1437 = s2_reg_dirty ? plru1_33 : _GEN_1244; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1438 = s2_reg_dirty ? plru1_34 : _GEN_1245; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1439 = s2_reg_dirty ? plru1_35 : _GEN_1246; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1440 = s2_reg_dirty ? plru1_36 : _GEN_1247; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1441 = s2_reg_dirty ? plru1_37 : _GEN_1248; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1442 = s2_reg_dirty ? plru1_38 : _GEN_1249; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1443 = s2_reg_dirty ? plru1_39 : _GEN_1250; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1444 = s2_reg_dirty ? plru1_40 : _GEN_1251; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1445 = s2_reg_dirty ? plru1_41 : _GEN_1252; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1446 = s2_reg_dirty ? plru1_42 : _GEN_1253; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1447 = s2_reg_dirty ? plru1_43 : _GEN_1254; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1448 = s2_reg_dirty ? plru1_44 : _GEN_1255; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1449 = s2_reg_dirty ? plru1_45 : _GEN_1256; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1450 = s2_reg_dirty ? plru1_46 : _GEN_1257; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1451 = s2_reg_dirty ? plru1_47 : _GEN_1258; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1452 = s2_reg_dirty ? plru1_48 : _GEN_1259; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1453 = s2_reg_dirty ? plru1_49 : _GEN_1260; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1454 = s2_reg_dirty ? plru1_50 : _GEN_1261; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1455 = s2_reg_dirty ? plru1_51 : _GEN_1262; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1456 = s2_reg_dirty ? plru1_52 : _GEN_1263; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1457 = s2_reg_dirty ? plru1_53 : _GEN_1264; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1458 = s2_reg_dirty ? plru1_54 : _GEN_1265; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1459 = s2_reg_dirty ? plru1_55 : _GEN_1266; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1460 = s2_reg_dirty ? plru1_56 : _GEN_1267; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1461 = s2_reg_dirty ? plru1_57 : _GEN_1268; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1462 = s2_reg_dirty ? plru1_58 : _GEN_1269; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1463 = s2_reg_dirty ? plru1_59 : _GEN_1270; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1464 = s2_reg_dirty ? plru1_60 : _GEN_1271; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1465 = s2_reg_dirty ? plru1_61 : _GEN_1272; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1466 = s2_reg_dirty ? plru1_62 : _GEN_1273; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1467 = s2_reg_dirty ? plru1_63 : _GEN_1274; // @[Cache.scala 349:27 Cache.scala 133:22]
  wire  _GEN_1468 = s2_reg_dirty ? plru2_0 : _GEN_1275; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1469 = s2_reg_dirty ? plru2_1 : _GEN_1276; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1470 = s2_reg_dirty ? plru2_2 : _GEN_1277; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1471 = s2_reg_dirty ? plru2_3 : _GEN_1278; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1472 = s2_reg_dirty ? plru2_4 : _GEN_1279; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1473 = s2_reg_dirty ? plru2_5 : _GEN_1280; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1474 = s2_reg_dirty ? plru2_6 : _GEN_1281; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1475 = s2_reg_dirty ? plru2_7 : _GEN_1282; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1476 = s2_reg_dirty ? plru2_8 : _GEN_1283; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1477 = s2_reg_dirty ? plru2_9 : _GEN_1284; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1478 = s2_reg_dirty ? plru2_10 : _GEN_1285; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1479 = s2_reg_dirty ? plru2_11 : _GEN_1286; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1480 = s2_reg_dirty ? plru2_12 : _GEN_1287; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1481 = s2_reg_dirty ? plru2_13 : _GEN_1288; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1482 = s2_reg_dirty ? plru2_14 : _GEN_1289; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1483 = s2_reg_dirty ? plru2_15 : _GEN_1290; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1484 = s2_reg_dirty ? plru2_16 : _GEN_1291; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1485 = s2_reg_dirty ? plru2_17 : _GEN_1292; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1486 = s2_reg_dirty ? plru2_18 : _GEN_1293; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1487 = s2_reg_dirty ? plru2_19 : _GEN_1294; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1488 = s2_reg_dirty ? plru2_20 : _GEN_1295; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1489 = s2_reg_dirty ? plru2_21 : _GEN_1296; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1490 = s2_reg_dirty ? plru2_22 : _GEN_1297; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1491 = s2_reg_dirty ? plru2_23 : _GEN_1298; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1492 = s2_reg_dirty ? plru2_24 : _GEN_1299; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1493 = s2_reg_dirty ? plru2_25 : _GEN_1300; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1494 = s2_reg_dirty ? plru2_26 : _GEN_1301; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1495 = s2_reg_dirty ? plru2_27 : _GEN_1302; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1496 = s2_reg_dirty ? plru2_28 : _GEN_1303; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1497 = s2_reg_dirty ? plru2_29 : _GEN_1304; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1498 = s2_reg_dirty ? plru2_30 : _GEN_1305; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1499 = s2_reg_dirty ? plru2_31 : _GEN_1306; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1500 = s2_reg_dirty ? plru2_32 : _GEN_1307; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1501 = s2_reg_dirty ? plru2_33 : _GEN_1308; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1502 = s2_reg_dirty ? plru2_34 : _GEN_1309; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1503 = s2_reg_dirty ? plru2_35 : _GEN_1310; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1504 = s2_reg_dirty ? plru2_36 : _GEN_1311; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1505 = s2_reg_dirty ? plru2_37 : _GEN_1312; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1506 = s2_reg_dirty ? plru2_38 : _GEN_1313; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1507 = s2_reg_dirty ? plru2_39 : _GEN_1314; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1508 = s2_reg_dirty ? plru2_40 : _GEN_1315; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1509 = s2_reg_dirty ? plru2_41 : _GEN_1316; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1510 = s2_reg_dirty ? plru2_42 : _GEN_1317; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1511 = s2_reg_dirty ? plru2_43 : _GEN_1318; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1512 = s2_reg_dirty ? plru2_44 : _GEN_1319; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1513 = s2_reg_dirty ? plru2_45 : _GEN_1320; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1514 = s2_reg_dirty ? plru2_46 : _GEN_1321; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1515 = s2_reg_dirty ? plru2_47 : _GEN_1322; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1516 = s2_reg_dirty ? plru2_48 : _GEN_1323; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1517 = s2_reg_dirty ? plru2_49 : _GEN_1324; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1518 = s2_reg_dirty ? plru2_50 : _GEN_1325; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1519 = s2_reg_dirty ? plru2_51 : _GEN_1326; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1520 = s2_reg_dirty ? plru2_52 : _GEN_1327; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1521 = s2_reg_dirty ? plru2_53 : _GEN_1328; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1522 = s2_reg_dirty ? plru2_54 : _GEN_1329; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1523 = s2_reg_dirty ? plru2_55 : _GEN_1330; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1524 = s2_reg_dirty ? plru2_56 : _GEN_1331; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1525 = s2_reg_dirty ? plru2_57 : _GEN_1332; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1526 = s2_reg_dirty ? plru2_58 : _GEN_1333; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1527 = s2_reg_dirty ? plru2_59 : _GEN_1334; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1528 = s2_reg_dirty ? plru2_60 : _GEN_1335; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1529 = s2_reg_dirty ? plru2_61 : _GEN_1336; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1530 = s2_reg_dirty ? plru2_62 : _GEN_1337; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _GEN_1531 = s2_reg_dirty ? plru2_63 : _GEN_1338; // @[Cache.scala 349:27 Cache.scala 135:22]
  wire  _T_23 = 4'h4 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_1532 = _T_12 ? 4'h5 : state; // @[Cache.scala 357:29 Cache.scala 358:15 Cache.scala 207:22]
  wire  _T_25 = 4'h5 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_1533 = _T_12 ? 4'h6 : state; // @[Cache.scala 362:29 Cache.scala 363:15 Cache.scala 207:22]
  wire  _T_27 = 4'h6 == state; // @[Conditional.scala 37:30]
  wire  _GEN_1854 = _T_14 ? _GEN_1019 : plru0_0; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1855 = _T_14 ? _GEN_1020 : plru0_1; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1856 = _T_14 ? _GEN_1021 : plru0_2; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1857 = _T_14 ? _GEN_1022 : plru0_3; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1858 = _T_14 ? _GEN_1023 : plru0_4; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1859 = _T_14 ? _GEN_1024 : plru0_5; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1860 = _T_14 ? _GEN_1025 : plru0_6; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1861 = _T_14 ? _GEN_1026 : plru0_7; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1862 = _T_14 ? _GEN_1027 : plru0_8; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1863 = _T_14 ? _GEN_1028 : plru0_9; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1864 = _T_14 ? _GEN_1029 : plru0_10; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1865 = _T_14 ? _GEN_1030 : plru0_11; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1866 = _T_14 ? _GEN_1031 : plru0_12; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1867 = _T_14 ? _GEN_1032 : plru0_13; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1868 = _T_14 ? _GEN_1033 : plru0_14; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1869 = _T_14 ? _GEN_1034 : plru0_15; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1870 = _T_14 ? _GEN_1035 : plru0_16; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1871 = _T_14 ? _GEN_1036 : plru0_17; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1872 = _T_14 ? _GEN_1037 : plru0_18; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1873 = _T_14 ? _GEN_1038 : plru0_19; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1874 = _T_14 ? _GEN_1039 : plru0_20; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1875 = _T_14 ? _GEN_1040 : plru0_21; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1876 = _T_14 ? _GEN_1041 : plru0_22; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1877 = _T_14 ? _GEN_1042 : plru0_23; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1878 = _T_14 ? _GEN_1043 : plru0_24; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1879 = _T_14 ? _GEN_1044 : plru0_25; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1880 = _T_14 ? _GEN_1045 : plru0_26; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1881 = _T_14 ? _GEN_1046 : plru0_27; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1882 = _T_14 ? _GEN_1047 : plru0_28; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1883 = _T_14 ? _GEN_1048 : plru0_29; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1884 = _T_14 ? _GEN_1049 : plru0_30; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1885 = _T_14 ? _GEN_1050 : plru0_31; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1886 = _T_14 ? _GEN_1051 : plru0_32; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1887 = _T_14 ? _GEN_1052 : plru0_33; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1888 = _T_14 ? _GEN_1053 : plru0_34; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1889 = _T_14 ? _GEN_1054 : plru0_35; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1890 = _T_14 ? _GEN_1055 : plru0_36; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1891 = _T_14 ? _GEN_1056 : plru0_37; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1892 = _T_14 ? _GEN_1057 : plru0_38; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1893 = _T_14 ? _GEN_1058 : plru0_39; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1894 = _T_14 ? _GEN_1059 : plru0_40; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1895 = _T_14 ? _GEN_1060 : plru0_41; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1896 = _T_14 ? _GEN_1061 : plru0_42; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1897 = _T_14 ? _GEN_1062 : plru0_43; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1898 = _T_14 ? _GEN_1063 : plru0_44; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1899 = _T_14 ? _GEN_1064 : plru0_45; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1900 = _T_14 ? _GEN_1065 : plru0_46; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1901 = _T_14 ? _GEN_1066 : plru0_47; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1902 = _T_14 ? _GEN_1067 : plru0_48; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1903 = _T_14 ? _GEN_1068 : plru0_49; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1904 = _T_14 ? _GEN_1069 : plru0_50; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1905 = _T_14 ? _GEN_1070 : plru0_51; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1906 = _T_14 ? _GEN_1071 : plru0_52; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1907 = _T_14 ? _GEN_1072 : plru0_53; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1908 = _T_14 ? _GEN_1073 : plru0_54; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1909 = _T_14 ? _GEN_1074 : plru0_55; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1910 = _T_14 ? _GEN_1075 : plru0_56; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1911 = _T_14 ? _GEN_1076 : plru0_57; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1912 = _T_14 ? _GEN_1077 : plru0_58; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1913 = _T_14 ? _GEN_1078 : plru0_59; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1914 = _T_14 ? _GEN_1079 : plru0_60; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1915 = _T_14 ? _GEN_1080 : plru0_61; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1916 = _T_14 ? _GEN_1081 : plru0_62; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1917 = _T_14 ? _GEN_1082 : plru0_63; // @[Cache.scala 368:30 Cache.scala 131:22]
  wire  _GEN_1918 = _T_14 ? _GEN_1211 : plru1_0; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1919 = _T_14 ? _GEN_1212 : plru1_1; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1920 = _T_14 ? _GEN_1213 : plru1_2; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1921 = _T_14 ? _GEN_1214 : plru1_3; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1922 = _T_14 ? _GEN_1215 : plru1_4; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1923 = _T_14 ? _GEN_1216 : plru1_5; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1924 = _T_14 ? _GEN_1217 : plru1_6; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1925 = _T_14 ? _GEN_1218 : plru1_7; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1926 = _T_14 ? _GEN_1219 : plru1_8; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1927 = _T_14 ? _GEN_1220 : plru1_9; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1928 = _T_14 ? _GEN_1221 : plru1_10; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1929 = _T_14 ? _GEN_1222 : plru1_11; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1930 = _T_14 ? _GEN_1223 : plru1_12; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1931 = _T_14 ? _GEN_1224 : plru1_13; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1932 = _T_14 ? _GEN_1225 : plru1_14; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1933 = _T_14 ? _GEN_1226 : plru1_15; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1934 = _T_14 ? _GEN_1227 : plru1_16; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1935 = _T_14 ? _GEN_1228 : plru1_17; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1936 = _T_14 ? _GEN_1229 : plru1_18; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1937 = _T_14 ? _GEN_1230 : plru1_19; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1938 = _T_14 ? _GEN_1231 : plru1_20; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1939 = _T_14 ? _GEN_1232 : plru1_21; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1940 = _T_14 ? _GEN_1233 : plru1_22; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1941 = _T_14 ? _GEN_1234 : plru1_23; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1942 = _T_14 ? _GEN_1235 : plru1_24; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1943 = _T_14 ? _GEN_1236 : plru1_25; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1944 = _T_14 ? _GEN_1237 : plru1_26; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1945 = _T_14 ? _GEN_1238 : plru1_27; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1946 = _T_14 ? _GEN_1239 : plru1_28; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1947 = _T_14 ? _GEN_1240 : plru1_29; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1948 = _T_14 ? _GEN_1241 : plru1_30; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1949 = _T_14 ? _GEN_1242 : plru1_31; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1950 = _T_14 ? _GEN_1243 : plru1_32; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1951 = _T_14 ? _GEN_1244 : plru1_33; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1952 = _T_14 ? _GEN_1245 : plru1_34; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1953 = _T_14 ? _GEN_1246 : plru1_35; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1954 = _T_14 ? _GEN_1247 : plru1_36; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1955 = _T_14 ? _GEN_1248 : plru1_37; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1956 = _T_14 ? _GEN_1249 : plru1_38; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1957 = _T_14 ? _GEN_1250 : plru1_39; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1958 = _T_14 ? _GEN_1251 : plru1_40; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1959 = _T_14 ? _GEN_1252 : plru1_41; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1960 = _T_14 ? _GEN_1253 : plru1_42; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1961 = _T_14 ? _GEN_1254 : plru1_43; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1962 = _T_14 ? _GEN_1255 : plru1_44; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1963 = _T_14 ? _GEN_1256 : plru1_45; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1964 = _T_14 ? _GEN_1257 : plru1_46; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1965 = _T_14 ? _GEN_1258 : plru1_47; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1966 = _T_14 ? _GEN_1259 : plru1_48; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1967 = _T_14 ? _GEN_1260 : plru1_49; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1968 = _T_14 ? _GEN_1261 : plru1_50; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1969 = _T_14 ? _GEN_1262 : plru1_51; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1970 = _T_14 ? _GEN_1263 : plru1_52; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1971 = _T_14 ? _GEN_1264 : plru1_53; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1972 = _T_14 ? _GEN_1265 : plru1_54; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1973 = _T_14 ? _GEN_1266 : plru1_55; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1974 = _T_14 ? _GEN_1267 : plru1_56; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1975 = _T_14 ? _GEN_1268 : plru1_57; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1976 = _T_14 ? _GEN_1269 : plru1_58; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1977 = _T_14 ? _GEN_1270 : plru1_59; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1978 = _T_14 ? _GEN_1271 : plru1_60; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1979 = _T_14 ? _GEN_1272 : plru1_61; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1980 = _T_14 ? _GEN_1273 : plru1_62; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1981 = _T_14 ? _GEN_1274 : plru1_63; // @[Cache.scala 368:30 Cache.scala 133:22]
  wire  _GEN_1982 = _T_14 ? _GEN_1275 : plru2_0; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1983 = _T_14 ? _GEN_1276 : plru2_1; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1984 = _T_14 ? _GEN_1277 : plru2_2; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1985 = _T_14 ? _GEN_1278 : plru2_3; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1986 = _T_14 ? _GEN_1279 : plru2_4; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1987 = _T_14 ? _GEN_1280 : plru2_5; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1988 = _T_14 ? _GEN_1281 : plru2_6; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1989 = _T_14 ? _GEN_1282 : plru2_7; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1990 = _T_14 ? _GEN_1283 : plru2_8; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1991 = _T_14 ? _GEN_1284 : plru2_9; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1992 = _T_14 ? _GEN_1285 : plru2_10; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1993 = _T_14 ? _GEN_1286 : plru2_11; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1994 = _T_14 ? _GEN_1287 : plru2_12; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1995 = _T_14 ? _GEN_1288 : plru2_13; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1996 = _T_14 ? _GEN_1289 : plru2_14; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1997 = _T_14 ? _GEN_1290 : plru2_15; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1998 = _T_14 ? _GEN_1291 : plru2_16; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_1999 = _T_14 ? _GEN_1292 : plru2_17; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2000 = _T_14 ? _GEN_1293 : plru2_18; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2001 = _T_14 ? _GEN_1294 : plru2_19; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2002 = _T_14 ? _GEN_1295 : plru2_20; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2003 = _T_14 ? _GEN_1296 : plru2_21; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2004 = _T_14 ? _GEN_1297 : plru2_22; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2005 = _T_14 ? _GEN_1298 : plru2_23; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2006 = _T_14 ? _GEN_1299 : plru2_24; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2007 = _T_14 ? _GEN_1300 : plru2_25; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2008 = _T_14 ? _GEN_1301 : plru2_26; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2009 = _T_14 ? _GEN_1302 : plru2_27; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2010 = _T_14 ? _GEN_1303 : plru2_28; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2011 = _T_14 ? _GEN_1304 : plru2_29; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2012 = _T_14 ? _GEN_1305 : plru2_30; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2013 = _T_14 ? _GEN_1306 : plru2_31; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2014 = _T_14 ? _GEN_1307 : plru2_32; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2015 = _T_14 ? _GEN_1308 : plru2_33; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2016 = _T_14 ? _GEN_1309 : plru2_34; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2017 = _T_14 ? _GEN_1310 : plru2_35; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2018 = _T_14 ? _GEN_1311 : plru2_36; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2019 = _T_14 ? _GEN_1312 : plru2_37; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2020 = _T_14 ? _GEN_1313 : plru2_38; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2021 = _T_14 ? _GEN_1314 : plru2_39; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2022 = _T_14 ? _GEN_1315 : plru2_40; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2023 = _T_14 ? _GEN_1316 : plru2_41; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2024 = _T_14 ? _GEN_1317 : plru2_42; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2025 = _T_14 ? _GEN_1318 : plru2_43; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2026 = _T_14 ? _GEN_1319 : plru2_44; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2027 = _T_14 ? _GEN_1320 : plru2_45; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2028 = _T_14 ? _GEN_1321 : plru2_46; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2029 = _T_14 ? _GEN_1322 : plru2_47; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2030 = _T_14 ? _GEN_1323 : plru2_48; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2031 = _T_14 ? _GEN_1324 : plru2_49; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2032 = _T_14 ? _GEN_1325 : plru2_50; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2033 = _T_14 ? _GEN_1326 : plru2_51; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2034 = _T_14 ? _GEN_1327 : plru2_52; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2035 = _T_14 ? _GEN_1328 : plru2_53; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2036 = _T_14 ? _GEN_1329 : plru2_54; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2037 = _T_14 ? _GEN_1330 : plru2_55; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2038 = _T_14 ? _GEN_1331 : plru2_56; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2039 = _T_14 ? _GEN_1332 : plru2_57; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2040 = _T_14 ? _GEN_1333 : plru2_58; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2041 = _T_14 ? _GEN_1334 : plru2_59; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2042 = _T_14 ? _GEN_1335 : plru2_60; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2043 = _T_14 ? _GEN_1336 : plru2_61; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2044 = _T_14 ? _GEN_1337 : plru2_62; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire  _GEN_2045 = _T_14 ? _GEN_1338 : plru2_63; // @[Cache.scala 368:30 Cache.scala 135:22]
  wire [3:0] _GEN_2046 = _T_14 ? 4'h7 : state; // @[Cache.scala 368:30 Cache.scala 370:15 Cache.scala 207:22]
  wire  _T_31 = 4'h7 == state; // @[Conditional.scala 37:30]
  reg [63:0] io_in_resp_bits_rdata_REG; // @[Cache.scala 374:36]
  wire  _T_32 = io_in_resp_ready & io_in_resp_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_2047 = _T_32 ? 4'h8 : state; // @[Cache.scala 375:29 Cache.scala 376:15 Cache.scala 207:22]
  wire [63:0] _GEN_2048 = _T_31 ? io_in_resp_bits_rdata_REG : 64'h0; // @[Conditional.scala 39:67 Cache.scala 374:26 Cache.scala 277:22]
  wire [3:0] _GEN_2049 = _T_31 ? _GEN_2047 : state; // @[Conditional.scala 39:67 Cache.scala 207:22]
  wire  _GEN_2050 = _T_27 ? 1'h0 : _GEN_27; // @[Conditional.scala 39:67 Cache.scala 367:14]
  wire  _GEN_2051 = _T_27 ? _GEN_1854 : plru0_0; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2052 = _T_27 ? _GEN_1855 : plru0_1; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2053 = _T_27 ? _GEN_1856 : plru0_2; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2054 = _T_27 ? _GEN_1857 : plru0_3; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2055 = _T_27 ? _GEN_1858 : plru0_4; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2056 = _T_27 ? _GEN_1859 : plru0_5; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2057 = _T_27 ? _GEN_1860 : plru0_6; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2058 = _T_27 ? _GEN_1861 : plru0_7; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2059 = _T_27 ? _GEN_1862 : plru0_8; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2060 = _T_27 ? _GEN_1863 : plru0_9; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2061 = _T_27 ? _GEN_1864 : plru0_10; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2062 = _T_27 ? _GEN_1865 : plru0_11; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2063 = _T_27 ? _GEN_1866 : plru0_12; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2064 = _T_27 ? _GEN_1867 : plru0_13; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2065 = _T_27 ? _GEN_1868 : plru0_14; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2066 = _T_27 ? _GEN_1869 : plru0_15; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2067 = _T_27 ? _GEN_1870 : plru0_16; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2068 = _T_27 ? _GEN_1871 : plru0_17; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2069 = _T_27 ? _GEN_1872 : plru0_18; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2070 = _T_27 ? _GEN_1873 : plru0_19; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2071 = _T_27 ? _GEN_1874 : plru0_20; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2072 = _T_27 ? _GEN_1875 : plru0_21; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2073 = _T_27 ? _GEN_1876 : plru0_22; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2074 = _T_27 ? _GEN_1877 : plru0_23; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2075 = _T_27 ? _GEN_1878 : plru0_24; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2076 = _T_27 ? _GEN_1879 : plru0_25; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2077 = _T_27 ? _GEN_1880 : plru0_26; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2078 = _T_27 ? _GEN_1881 : plru0_27; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2079 = _T_27 ? _GEN_1882 : plru0_28; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2080 = _T_27 ? _GEN_1883 : plru0_29; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2081 = _T_27 ? _GEN_1884 : plru0_30; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2082 = _T_27 ? _GEN_1885 : plru0_31; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2083 = _T_27 ? _GEN_1886 : plru0_32; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2084 = _T_27 ? _GEN_1887 : plru0_33; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2085 = _T_27 ? _GEN_1888 : plru0_34; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2086 = _T_27 ? _GEN_1889 : plru0_35; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2087 = _T_27 ? _GEN_1890 : plru0_36; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2088 = _T_27 ? _GEN_1891 : plru0_37; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2089 = _T_27 ? _GEN_1892 : plru0_38; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2090 = _T_27 ? _GEN_1893 : plru0_39; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2091 = _T_27 ? _GEN_1894 : plru0_40; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2092 = _T_27 ? _GEN_1895 : plru0_41; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2093 = _T_27 ? _GEN_1896 : plru0_42; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2094 = _T_27 ? _GEN_1897 : plru0_43; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2095 = _T_27 ? _GEN_1898 : plru0_44; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2096 = _T_27 ? _GEN_1899 : plru0_45; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2097 = _T_27 ? _GEN_1900 : plru0_46; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2098 = _T_27 ? _GEN_1901 : plru0_47; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2099 = _T_27 ? _GEN_1902 : plru0_48; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2100 = _T_27 ? _GEN_1903 : plru0_49; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2101 = _T_27 ? _GEN_1904 : plru0_50; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2102 = _T_27 ? _GEN_1905 : plru0_51; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2103 = _T_27 ? _GEN_1906 : plru0_52; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2104 = _T_27 ? _GEN_1907 : plru0_53; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2105 = _T_27 ? _GEN_1908 : plru0_54; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2106 = _T_27 ? _GEN_1909 : plru0_55; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2107 = _T_27 ? _GEN_1910 : plru0_56; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2108 = _T_27 ? _GEN_1911 : plru0_57; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2109 = _T_27 ? _GEN_1912 : plru0_58; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2110 = _T_27 ? _GEN_1913 : plru0_59; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2111 = _T_27 ? _GEN_1914 : plru0_60; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2112 = _T_27 ? _GEN_1915 : plru0_61; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2113 = _T_27 ? _GEN_1916 : plru0_62; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2114 = _T_27 ? _GEN_1917 : plru0_63; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2115 = _T_27 ? _GEN_1918 : plru1_0; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2116 = _T_27 ? _GEN_1919 : plru1_1; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2117 = _T_27 ? _GEN_1920 : plru1_2; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2118 = _T_27 ? _GEN_1921 : plru1_3; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2119 = _T_27 ? _GEN_1922 : plru1_4; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2120 = _T_27 ? _GEN_1923 : plru1_5; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2121 = _T_27 ? _GEN_1924 : plru1_6; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2122 = _T_27 ? _GEN_1925 : plru1_7; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2123 = _T_27 ? _GEN_1926 : plru1_8; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2124 = _T_27 ? _GEN_1927 : plru1_9; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2125 = _T_27 ? _GEN_1928 : plru1_10; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2126 = _T_27 ? _GEN_1929 : plru1_11; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2127 = _T_27 ? _GEN_1930 : plru1_12; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2128 = _T_27 ? _GEN_1931 : plru1_13; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2129 = _T_27 ? _GEN_1932 : plru1_14; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2130 = _T_27 ? _GEN_1933 : plru1_15; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2131 = _T_27 ? _GEN_1934 : plru1_16; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2132 = _T_27 ? _GEN_1935 : plru1_17; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2133 = _T_27 ? _GEN_1936 : plru1_18; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2134 = _T_27 ? _GEN_1937 : plru1_19; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2135 = _T_27 ? _GEN_1938 : plru1_20; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2136 = _T_27 ? _GEN_1939 : plru1_21; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2137 = _T_27 ? _GEN_1940 : plru1_22; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2138 = _T_27 ? _GEN_1941 : plru1_23; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2139 = _T_27 ? _GEN_1942 : plru1_24; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2140 = _T_27 ? _GEN_1943 : plru1_25; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2141 = _T_27 ? _GEN_1944 : plru1_26; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2142 = _T_27 ? _GEN_1945 : plru1_27; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2143 = _T_27 ? _GEN_1946 : plru1_28; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2144 = _T_27 ? _GEN_1947 : plru1_29; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2145 = _T_27 ? _GEN_1948 : plru1_30; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2146 = _T_27 ? _GEN_1949 : plru1_31; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2147 = _T_27 ? _GEN_1950 : plru1_32; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2148 = _T_27 ? _GEN_1951 : plru1_33; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2149 = _T_27 ? _GEN_1952 : plru1_34; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2150 = _T_27 ? _GEN_1953 : plru1_35; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2151 = _T_27 ? _GEN_1954 : plru1_36; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2152 = _T_27 ? _GEN_1955 : plru1_37; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2153 = _T_27 ? _GEN_1956 : plru1_38; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2154 = _T_27 ? _GEN_1957 : plru1_39; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2155 = _T_27 ? _GEN_1958 : plru1_40; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2156 = _T_27 ? _GEN_1959 : plru1_41; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2157 = _T_27 ? _GEN_1960 : plru1_42; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2158 = _T_27 ? _GEN_1961 : plru1_43; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2159 = _T_27 ? _GEN_1962 : plru1_44; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2160 = _T_27 ? _GEN_1963 : plru1_45; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2161 = _T_27 ? _GEN_1964 : plru1_46; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2162 = _T_27 ? _GEN_1965 : plru1_47; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2163 = _T_27 ? _GEN_1966 : plru1_48; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2164 = _T_27 ? _GEN_1967 : plru1_49; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2165 = _T_27 ? _GEN_1968 : plru1_50; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2166 = _T_27 ? _GEN_1969 : plru1_51; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2167 = _T_27 ? _GEN_1970 : plru1_52; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2168 = _T_27 ? _GEN_1971 : plru1_53; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2169 = _T_27 ? _GEN_1972 : plru1_54; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2170 = _T_27 ? _GEN_1973 : plru1_55; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2171 = _T_27 ? _GEN_1974 : plru1_56; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2172 = _T_27 ? _GEN_1975 : plru1_57; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2173 = _T_27 ? _GEN_1976 : plru1_58; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2174 = _T_27 ? _GEN_1977 : plru1_59; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2175 = _T_27 ? _GEN_1978 : plru1_60; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2176 = _T_27 ? _GEN_1979 : plru1_61; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2177 = _T_27 ? _GEN_1980 : plru1_62; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2178 = _T_27 ? _GEN_1981 : plru1_63; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2179 = _T_27 ? _GEN_1982 : plru2_0; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2180 = _T_27 ? _GEN_1983 : plru2_1; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2181 = _T_27 ? _GEN_1984 : plru2_2; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2182 = _T_27 ? _GEN_1985 : plru2_3; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2183 = _T_27 ? _GEN_1986 : plru2_4; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2184 = _T_27 ? _GEN_1987 : plru2_5; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2185 = _T_27 ? _GEN_1988 : plru2_6; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2186 = _T_27 ? _GEN_1989 : plru2_7; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2187 = _T_27 ? _GEN_1990 : plru2_8; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2188 = _T_27 ? _GEN_1991 : plru2_9; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2189 = _T_27 ? _GEN_1992 : plru2_10; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2190 = _T_27 ? _GEN_1993 : plru2_11; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2191 = _T_27 ? _GEN_1994 : plru2_12; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2192 = _T_27 ? _GEN_1995 : plru2_13; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2193 = _T_27 ? _GEN_1996 : plru2_14; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2194 = _T_27 ? _GEN_1997 : plru2_15; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2195 = _T_27 ? _GEN_1998 : plru2_16; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2196 = _T_27 ? _GEN_1999 : plru2_17; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2197 = _T_27 ? _GEN_2000 : plru2_18; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2198 = _T_27 ? _GEN_2001 : plru2_19; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2199 = _T_27 ? _GEN_2002 : plru2_20; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2200 = _T_27 ? _GEN_2003 : plru2_21; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2201 = _T_27 ? _GEN_2004 : plru2_22; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2202 = _T_27 ? _GEN_2005 : plru2_23; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2203 = _T_27 ? _GEN_2006 : plru2_24; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2204 = _T_27 ? _GEN_2007 : plru2_25; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2205 = _T_27 ? _GEN_2008 : plru2_26; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2206 = _T_27 ? _GEN_2009 : plru2_27; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2207 = _T_27 ? _GEN_2010 : plru2_28; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2208 = _T_27 ? _GEN_2011 : plru2_29; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2209 = _T_27 ? _GEN_2012 : plru2_30; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2210 = _T_27 ? _GEN_2013 : plru2_31; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2211 = _T_27 ? _GEN_2014 : plru2_32; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2212 = _T_27 ? _GEN_2015 : plru2_33; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2213 = _T_27 ? _GEN_2016 : plru2_34; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2214 = _T_27 ? _GEN_2017 : plru2_35; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2215 = _T_27 ? _GEN_2018 : plru2_36; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2216 = _T_27 ? _GEN_2019 : plru2_37; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2217 = _T_27 ? _GEN_2020 : plru2_38; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2218 = _T_27 ? _GEN_2021 : plru2_39; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2219 = _T_27 ? _GEN_2022 : plru2_40; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2220 = _T_27 ? _GEN_2023 : plru2_41; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2221 = _T_27 ? _GEN_2024 : plru2_42; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2222 = _T_27 ? _GEN_2025 : plru2_43; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2223 = _T_27 ? _GEN_2026 : plru2_44; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2224 = _T_27 ? _GEN_2027 : plru2_45; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2225 = _T_27 ? _GEN_2028 : plru2_46; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2226 = _T_27 ? _GEN_2029 : plru2_47; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2227 = _T_27 ? _GEN_2030 : plru2_48; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2228 = _T_27 ? _GEN_2031 : plru2_49; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2229 = _T_27 ? _GEN_2032 : plru2_50; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2230 = _T_27 ? _GEN_2033 : plru2_51; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2231 = _T_27 ? _GEN_2034 : plru2_52; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2232 = _T_27 ? _GEN_2035 : plru2_53; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2233 = _T_27 ? _GEN_2036 : plru2_54; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2234 = _T_27 ? _GEN_2037 : plru2_55; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2235 = _T_27 ? _GEN_2038 : plru2_56; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2236 = _T_27 ? _GEN_2039 : plru2_57; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2237 = _T_27 ? _GEN_2040 : plru2_58; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2238 = _T_27 ? _GEN_2041 : plru2_59; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2239 = _T_27 ? _GEN_2042 : plru2_60; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2240 = _T_27 ? _GEN_2043 : plru2_61; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2241 = _T_27 ? _GEN_2044 : plru2_62; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2242 = _T_27 ? _GEN_2045 : plru2_63; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire [3:0] _GEN_2243 = _T_27 ? _GEN_2046 : _GEN_2049; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_2244 = _T_27 ? 64'h0 : _GEN_2048; // @[Conditional.scala 39:67 Cache.scala 277:22]
  wire [3:0] _GEN_2245 = _T_25 ? _GEN_1533 : _GEN_2243; // @[Conditional.scala 39:67]
  wire  _GEN_2246 = _T_25 ? _GEN_27 : _GEN_2050; // @[Conditional.scala 39:67]
  wire  _GEN_2247 = _T_25 ? plru0_0 : _GEN_2051; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2248 = _T_25 ? plru0_1 : _GEN_2052; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2249 = _T_25 ? plru0_2 : _GEN_2053; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2250 = _T_25 ? plru0_3 : _GEN_2054; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2251 = _T_25 ? plru0_4 : _GEN_2055; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2252 = _T_25 ? plru0_5 : _GEN_2056; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2253 = _T_25 ? plru0_6 : _GEN_2057; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2254 = _T_25 ? plru0_7 : _GEN_2058; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2255 = _T_25 ? plru0_8 : _GEN_2059; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2256 = _T_25 ? plru0_9 : _GEN_2060; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2257 = _T_25 ? plru0_10 : _GEN_2061; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2258 = _T_25 ? plru0_11 : _GEN_2062; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2259 = _T_25 ? plru0_12 : _GEN_2063; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2260 = _T_25 ? plru0_13 : _GEN_2064; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2261 = _T_25 ? plru0_14 : _GEN_2065; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2262 = _T_25 ? plru0_15 : _GEN_2066; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2263 = _T_25 ? plru0_16 : _GEN_2067; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2264 = _T_25 ? plru0_17 : _GEN_2068; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2265 = _T_25 ? plru0_18 : _GEN_2069; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2266 = _T_25 ? plru0_19 : _GEN_2070; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2267 = _T_25 ? plru0_20 : _GEN_2071; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2268 = _T_25 ? plru0_21 : _GEN_2072; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2269 = _T_25 ? plru0_22 : _GEN_2073; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2270 = _T_25 ? plru0_23 : _GEN_2074; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2271 = _T_25 ? plru0_24 : _GEN_2075; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2272 = _T_25 ? plru0_25 : _GEN_2076; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2273 = _T_25 ? plru0_26 : _GEN_2077; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2274 = _T_25 ? plru0_27 : _GEN_2078; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2275 = _T_25 ? plru0_28 : _GEN_2079; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2276 = _T_25 ? plru0_29 : _GEN_2080; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2277 = _T_25 ? plru0_30 : _GEN_2081; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2278 = _T_25 ? plru0_31 : _GEN_2082; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2279 = _T_25 ? plru0_32 : _GEN_2083; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2280 = _T_25 ? plru0_33 : _GEN_2084; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2281 = _T_25 ? plru0_34 : _GEN_2085; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2282 = _T_25 ? plru0_35 : _GEN_2086; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2283 = _T_25 ? plru0_36 : _GEN_2087; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2284 = _T_25 ? plru0_37 : _GEN_2088; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2285 = _T_25 ? plru0_38 : _GEN_2089; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2286 = _T_25 ? plru0_39 : _GEN_2090; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2287 = _T_25 ? plru0_40 : _GEN_2091; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2288 = _T_25 ? plru0_41 : _GEN_2092; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2289 = _T_25 ? plru0_42 : _GEN_2093; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2290 = _T_25 ? plru0_43 : _GEN_2094; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2291 = _T_25 ? plru0_44 : _GEN_2095; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2292 = _T_25 ? plru0_45 : _GEN_2096; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2293 = _T_25 ? plru0_46 : _GEN_2097; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2294 = _T_25 ? plru0_47 : _GEN_2098; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2295 = _T_25 ? plru0_48 : _GEN_2099; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2296 = _T_25 ? plru0_49 : _GEN_2100; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2297 = _T_25 ? plru0_50 : _GEN_2101; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2298 = _T_25 ? plru0_51 : _GEN_2102; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2299 = _T_25 ? plru0_52 : _GEN_2103; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2300 = _T_25 ? plru0_53 : _GEN_2104; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2301 = _T_25 ? plru0_54 : _GEN_2105; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2302 = _T_25 ? plru0_55 : _GEN_2106; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2303 = _T_25 ? plru0_56 : _GEN_2107; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2304 = _T_25 ? plru0_57 : _GEN_2108; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2305 = _T_25 ? plru0_58 : _GEN_2109; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2306 = _T_25 ? plru0_59 : _GEN_2110; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2307 = _T_25 ? plru0_60 : _GEN_2111; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2308 = _T_25 ? plru0_61 : _GEN_2112; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2309 = _T_25 ? plru0_62 : _GEN_2113; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2310 = _T_25 ? plru0_63 : _GEN_2114; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2311 = _T_25 ? plru1_0 : _GEN_2115; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2312 = _T_25 ? plru1_1 : _GEN_2116; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2313 = _T_25 ? plru1_2 : _GEN_2117; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2314 = _T_25 ? plru1_3 : _GEN_2118; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2315 = _T_25 ? plru1_4 : _GEN_2119; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2316 = _T_25 ? plru1_5 : _GEN_2120; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2317 = _T_25 ? plru1_6 : _GEN_2121; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2318 = _T_25 ? plru1_7 : _GEN_2122; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2319 = _T_25 ? plru1_8 : _GEN_2123; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2320 = _T_25 ? plru1_9 : _GEN_2124; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2321 = _T_25 ? plru1_10 : _GEN_2125; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2322 = _T_25 ? plru1_11 : _GEN_2126; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2323 = _T_25 ? plru1_12 : _GEN_2127; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2324 = _T_25 ? plru1_13 : _GEN_2128; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2325 = _T_25 ? plru1_14 : _GEN_2129; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2326 = _T_25 ? plru1_15 : _GEN_2130; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2327 = _T_25 ? plru1_16 : _GEN_2131; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2328 = _T_25 ? plru1_17 : _GEN_2132; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2329 = _T_25 ? plru1_18 : _GEN_2133; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2330 = _T_25 ? plru1_19 : _GEN_2134; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2331 = _T_25 ? plru1_20 : _GEN_2135; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2332 = _T_25 ? plru1_21 : _GEN_2136; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2333 = _T_25 ? plru1_22 : _GEN_2137; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2334 = _T_25 ? plru1_23 : _GEN_2138; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2335 = _T_25 ? plru1_24 : _GEN_2139; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2336 = _T_25 ? plru1_25 : _GEN_2140; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2337 = _T_25 ? plru1_26 : _GEN_2141; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2338 = _T_25 ? plru1_27 : _GEN_2142; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2339 = _T_25 ? plru1_28 : _GEN_2143; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2340 = _T_25 ? plru1_29 : _GEN_2144; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2341 = _T_25 ? plru1_30 : _GEN_2145; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2342 = _T_25 ? plru1_31 : _GEN_2146; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2343 = _T_25 ? plru1_32 : _GEN_2147; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2344 = _T_25 ? plru1_33 : _GEN_2148; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2345 = _T_25 ? plru1_34 : _GEN_2149; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2346 = _T_25 ? plru1_35 : _GEN_2150; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2347 = _T_25 ? plru1_36 : _GEN_2151; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2348 = _T_25 ? plru1_37 : _GEN_2152; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2349 = _T_25 ? plru1_38 : _GEN_2153; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2350 = _T_25 ? plru1_39 : _GEN_2154; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2351 = _T_25 ? plru1_40 : _GEN_2155; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2352 = _T_25 ? plru1_41 : _GEN_2156; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2353 = _T_25 ? plru1_42 : _GEN_2157; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2354 = _T_25 ? plru1_43 : _GEN_2158; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2355 = _T_25 ? plru1_44 : _GEN_2159; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2356 = _T_25 ? plru1_45 : _GEN_2160; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2357 = _T_25 ? plru1_46 : _GEN_2161; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2358 = _T_25 ? plru1_47 : _GEN_2162; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2359 = _T_25 ? plru1_48 : _GEN_2163; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2360 = _T_25 ? plru1_49 : _GEN_2164; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2361 = _T_25 ? plru1_50 : _GEN_2165; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2362 = _T_25 ? plru1_51 : _GEN_2166; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2363 = _T_25 ? plru1_52 : _GEN_2167; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2364 = _T_25 ? plru1_53 : _GEN_2168; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2365 = _T_25 ? plru1_54 : _GEN_2169; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2366 = _T_25 ? plru1_55 : _GEN_2170; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2367 = _T_25 ? plru1_56 : _GEN_2171; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2368 = _T_25 ? plru1_57 : _GEN_2172; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2369 = _T_25 ? plru1_58 : _GEN_2173; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2370 = _T_25 ? plru1_59 : _GEN_2174; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2371 = _T_25 ? plru1_60 : _GEN_2175; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2372 = _T_25 ? plru1_61 : _GEN_2176; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2373 = _T_25 ? plru1_62 : _GEN_2177; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2374 = _T_25 ? plru1_63 : _GEN_2178; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2375 = _T_25 ? plru2_0 : _GEN_2179; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2376 = _T_25 ? plru2_1 : _GEN_2180; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2377 = _T_25 ? plru2_2 : _GEN_2181; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2378 = _T_25 ? plru2_3 : _GEN_2182; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2379 = _T_25 ? plru2_4 : _GEN_2183; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2380 = _T_25 ? plru2_5 : _GEN_2184; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2381 = _T_25 ? plru2_6 : _GEN_2185; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2382 = _T_25 ? plru2_7 : _GEN_2186; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2383 = _T_25 ? plru2_8 : _GEN_2187; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2384 = _T_25 ? plru2_9 : _GEN_2188; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2385 = _T_25 ? plru2_10 : _GEN_2189; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2386 = _T_25 ? plru2_11 : _GEN_2190; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2387 = _T_25 ? plru2_12 : _GEN_2191; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2388 = _T_25 ? plru2_13 : _GEN_2192; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2389 = _T_25 ? plru2_14 : _GEN_2193; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2390 = _T_25 ? plru2_15 : _GEN_2194; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2391 = _T_25 ? plru2_16 : _GEN_2195; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2392 = _T_25 ? plru2_17 : _GEN_2196; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2393 = _T_25 ? plru2_18 : _GEN_2197; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2394 = _T_25 ? plru2_19 : _GEN_2198; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2395 = _T_25 ? plru2_20 : _GEN_2199; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2396 = _T_25 ? plru2_21 : _GEN_2200; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2397 = _T_25 ? plru2_22 : _GEN_2201; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2398 = _T_25 ? plru2_23 : _GEN_2202; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2399 = _T_25 ? plru2_24 : _GEN_2203; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2400 = _T_25 ? plru2_25 : _GEN_2204; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2401 = _T_25 ? plru2_26 : _GEN_2205; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2402 = _T_25 ? plru2_27 : _GEN_2206; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2403 = _T_25 ? plru2_28 : _GEN_2207; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2404 = _T_25 ? plru2_29 : _GEN_2208; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2405 = _T_25 ? plru2_30 : _GEN_2209; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2406 = _T_25 ? plru2_31 : _GEN_2210; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2407 = _T_25 ? plru2_32 : _GEN_2211; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2408 = _T_25 ? plru2_33 : _GEN_2212; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2409 = _T_25 ? plru2_34 : _GEN_2213; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2410 = _T_25 ? plru2_35 : _GEN_2214; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2411 = _T_25 ? plru2_36 : _GEN_2215; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2412 = _T_25 ? plru2_37 : _GEN_2216; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2413 = _T_25 ? plru2_38 : _GEN_2217; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2414 = _T_25 ? plru2_39 : _GEN_2218; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2415 = _T_25 ? plru2_40 : _GEN_2219; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2416 = _T_25 ? plru2_41 : _GEN_2220; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2417 = _T_25 ? plru2_42 : _GEN_2221; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2418 = _T_25 ? plru2_43 : _GEN_2222; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2419 = _T_25 ? plru2_44 : _GEN_2223; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2420 = _T_25 ? plru2_45 : _GEN_2224; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2421 = _T_25 ? plru2_46 : _GEN_2225; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2422 = _T_25 ? plru2_47 : _GEN_2226; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2423 = _T_25 ? plru2_48 : _GEN_2227; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2424 = _T_25 ? plru2_49 : _GEN_2228; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2425 = _T_25 ? plru2_50 : _GEN_2229; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2426 = _T_25 ? plru2_51 : _GEN_2230; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2427 = _T_25 ? plru2_52 : _GEN_2231; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2428 = _T_25 ? plru2_53 : _GEN_2232; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2429 = _T_25 ? plru2_54 : _GEN_2233; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2430 = _T_25 ? plru2_55 : _GEN_2234; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2431 = _T_25 ? plru2_56 : _GEN_2235; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2432 = _T_25 ? plru2_57 : _GEN_2236; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2433 = _T_25 ? plru2_58 : _GEN_2237; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2434 = _T_25 ? plru2_59 : _GEN_2238; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2435 = _T_25 ? plru2_60 : _GEN_2239; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2436 = _T_25 ? plru2_61 : _GEN_2240; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2437 = _T_25 ? plru2_62 : _GEN_2241; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2438 = _T_25 ? plru2_63 : _GEN_2242; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire [63:0] _GEN_2439 = _T_25 ? 64'h0 : _GEN_2244; // @[Conditional.scala 39:67 Cache.scala 277:22]
  wire [3:0] _GEN_2440 = _T_23 ? _GEN_1532 : _GEN_2245; // @[Conditional.scala 39:67]
  wire  _GEN_2441 = _T_23 ? _GEN_27 : _GEN_2246; // @[Conditional.scala 39:67]
  wire  _GEN_2442 = _T_23 ? plru0_0 : _GEN_2247; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2443 = _T_23 ? plru0_1 : _GEN_2248; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2444 = _T_23 ? plru0_2 : _GEN_2249; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2445 = _T_23 ? plru0_3 : _GEN_2250; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2446 = _T_23 ? plru0_4 : _GEN_2251; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2447 = _T_23 ? plru0_5 : _GEN_2252; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2448 = _T_23 ? plru0_6 : _GEN_2253; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2449 = _T_23 ? plru0_7 : _GEN_2254; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2450 = _T_23 ? plru0_8 : _GEN_2255; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2451 = _T_23 ? plru0_9 : _GEN_2256; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2452 = _T_23 ? plru0_10 : _GEN_2257; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2453 = _T_23 ? plru0_11 : _GEN_2258; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2454 = _T_23 ? plru0_12 : _GEN_2259; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2455 = _T_23 ? plru0_13 : _GEN_2260; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2456 = _T_23 ? plru0_14 : _GEN_2261; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2457 = _T_23 ? plru0_15 : _GEN_2262; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2458 = _T_23 ? plru0_16 : _GEN_2263; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2459 = _T_23 ? plru0_17 : _GEN_2264; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2460 = _T_23 ? plru0_18 : _GEN_2265; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2461 = _T_23 ? plru0_19 : _GEN_2266; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2462 = _T_23 ? plru0_20 : _GEN_2267; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2463 = _T_23 ? plru0_21 : _GEN_2268; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2464 = _T_23 ? plru0_22 : _GEN_2269; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2465 = _T_23 ? plru0_23 : _GEN_2270; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2466 = _T_23 ? plru0_24 : _GEN_2271; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2467 = _T_23 ? plru0_25 : _GEN_2272; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2468 = _T_23 ? plru0_26 : _GEN_2273; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2469 = _T_23 ? plru0_27 : _GEN_2274; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2470 = _T_23 ? plru0_28 : _GEN_2275; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2471 = _T_23 ? plru0_29 : _GEN_2276; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2472 = _T_23 ? plru0_30 : _GEN_2277; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2473 = _T_23 ? plru0_31 : _GEN_2278; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2474 = _T_23 ? plru0_32 : _GEN_2279; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2475 = _T_23 ? plru0_33 : _GEN_2280; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2476 = _T_23 ? plru0_34 : _GEN_2281; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2477 = _T_23 ? plru0_35 : _GEN_2282; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2478 = _T_23 ? plru0_36 : _GEN_2283; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2479 = _T_23 ? plru0_37 : _GEN_2284; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2480 = _T_23 ? plru0_38 : _GEN_2285; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2481 = _T_23 ? plru0_39 : _GEN_2286; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2482 = _T_23 ? plru0_40 : _GEN_2287; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2483 = _T_23 ? plru0_41 : _GEN_2288; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2484 = _T_23 ? plru0_42 : _GEN_2289; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2485 = _T_23 ? plru0_43 : _GEN_2290; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2486 = _T_23 ? plru0_44 : _GEN_2291; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2487 = _T_23 ? plru0_45 : _GEN_2292; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2488 = _T_23 ? plru0_46 : _GEN_2293; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2489 = _T_23 ? plru0_47 : _GEN_2294; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2490 = _T_23 ? plru0_48 : _GEN_2295; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2491 = _T_23 ? plru0_49 : _GEN_2296; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2492 = _T_23 ? plru0_50 : _GEN_2297; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2493 = _T_23 ? plru0_51 : _GEN_2298; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2494 = _T_23 ? plru0_52 : _GEN_2299; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2495 = _T_23 ? plru0_53 : _GEN_2300; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2496 = _T_23 ? plru0_54 : _GEN_2301; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2497 = _T_23 ? plru0_55 : _GEN_2302; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2498 = _T_23 ? plru0_56 : _GEN_2303; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2499 = _T_23 ? plru0_57 : _GEN_2304; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2500 = _T_23 ? plru0_58 : _GEN_2305; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2501 = _T_23 ? plru0_59 : _GEN_2306; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2502 = _T_23 ? plru0_60 : _GEN_2307; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2503 = _T_23 ? plru0_61 : _GEN_2308; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2504 = _T_23 ? plru0_62 : _GEN_2309; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2505 = _T_23 ? plru0_63 : _GEN_2310; // @[Conditional.scala 39:67 Cache.scala 131:22]
  wire  _GEN_2506 = _T_23 ? plru1_0 : _GEN_2311; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2507 = _T_23 ? plru1_1 : _GEN_2312; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2508 = _T_23 ? plru1_2 : _GEN_2313; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2509 = _T_23 ? plru1_3 : _GEN_2314; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2510 = _T_23 ? plru1_4 : _GEN_2315; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2511 = _T_23 ? plru1_5 : _GEN_2316; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2512 = _T_23 ? plru1_6 : _GEN_2317; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2513 = _T_23 ? plru1_7 : _GEN_2318; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2514 = _T_23 ? plru1_8 : _GEN_2319; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2515 = _T_23 ? plru1_9 : _GEN_2320; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2516 = _T_23 ? plru1_10 : _GEN_2321; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2517 = _T_23 ? plru1_11 : _GEN_2322; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2518 = _T_23 ? plru1_12 : _GEN_2323; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2519 = _T_23 ? plru1_13 : _GEN_2324; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2520 = _T_23 ? plru1_14 : _GEN_2325; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2521 = _T_23 ? plru1_15 : _GEN_2326; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2522 = _T_23 ? plru1_16 : _GEN_2327; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2523 = _T_23 ? plru1_17 : _GEN_2328; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2524 = _T_23 ? plru1_18 : _GEN_2329; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2525 = _T_23 ? plru1_19 : _GEN_2330; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2526 = _T_23 ? plru1_20 : _GEN_2331; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2527 = _T_23 ? plru1_21 : _GEN_2332; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2528 = _T_23 ? plru1_22 : _GEN_2333; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2529 = _T_23 ? plru1_23 : _GEN_2334; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2530 = _T_23 ? plru1_24 : _GEN_2335; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2531 = _T_23 ? plru1_25 : _GEN_2336; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2532 = _T_23 ? plru1_26 : _GEN_2337; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2533 = _T_23 ? plru1_27 : _GEN_2338; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2534 = _T_23 ? plru1_28 : _GEN_2339; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2535 = _T_23 ? plru1_29 : _GEN_2340; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2536 = _T_23 ? plru1_30 : _GEN_2341; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2537 = _T_23 ? plru1_31 : _GEN_2342; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2538 = _T_23 ? plru1_32 : _GEN_2343; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2539 = _T_23 ? plru1_33 : _GEN_2344; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2540 = _T_23 ? plru1_34 : _GEN_2345; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2541 = _T_23 ? plru1_35 : _GEN_2346; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2542 = _T_23 ? plru1_36 : _GEN_2347; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2543 = _T_23 ? plru1_37 : _GEN_2348; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2544 = _T_23 ? plru1_38 : _GEN_2349; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2545 = _T_23 ? plru1_39 : _GEN_2350; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2546 = _T_23 ? plru1_40 : _GEN_2351; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2547 = _T_23 ? plru1_41 : _GEN_2352; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2548 = _T_23 ? plru1_42 : _GEN_2353; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2549 = _T_23 ? plru1_43 : _GEN_2354; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2550 = _T_23 ? plru1_44 : _GEN_2355; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2551 = _T_23 ? plru1_45 : _GEN_2356; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2552 = _T_23 ? plru1_46 : _GEN_2357; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2553 = _T_23 ? plru1_47 : _GEN_2358; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2554 = _T_23 ? plru1_48 : _GEN_2359; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2555 = _T_23 ? plru1_49 : _GEN_2360; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2556 = _T_23 ? plru1_50 : _GEN_2361; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2557 = _T_23 ? plru1_51 : _GEN_2362; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2558 = _T_23 ? plru1_52 : _GEN_2363; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2559 = _T_23 ? plru1_53 : _GEN_2364; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2560 = _T_23 ? plru1_54 : _GEN_2365; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2561 = _T_23 ? plru1_55 : _GEN_2366; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2562 = _T_23 ? plru1_56 : _GEN_2367; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2563 = _T_23 ? plru1_57 : _GEN_2368; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2564 = _T_23 ? plru1_58 : _GEN_2369; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2565 = _T_23 ? plru1_59 : _GEN_2370; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2566 = _T_23 ? plru1_60 : _GEN_2371; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2567 = _T_23 ? plru1_61 : _GEN_2372; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2568 = _T_23 ? plru1_62 : _GEN_2373; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2569 = _T_23 ? plru1_63 : _GEN_2374; // @[Conditional.scala 39:67 Cache.scala 133:22]
  wire  _GEN_2570 = _T_23 ? plru2_0 : _GEN_2375; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2571 = _T_23 ? plru2_1 : _GEN_2376; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2572 = _T_23 ? plru2_2 : _GEN_2377; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2573 = _T_23 ? plru2_3 : _GEN_2378; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2574 = _T_23 ? plru2_4 : _GEN_2379; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2575 = _T_23 ? plru2_5 : _GEN_2380; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2576 = _T_23 ? plru2_6 : _GEN_2381; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2577 = _T_23 ? plru2_7 : _GEN_2382; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2578 = _T_23 ? plru2_8 : _GEN_2383; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2579 = _T_23 ? plru2_9 : _GEN_2384; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2580 = _T_23 ? plru2_10 : _GEN_2385; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2581 = _T_23 ? plru2_11 : _GEN_2386; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2582 = _T_23 ? plru2_12 : _GEN_2387; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2583 = _T_23 ? plru2_13 : _GEN_2388; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2584 = _T_23 ? plru2_14 : _GEN_2389; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2585 = _T_23 ? plru2_15 : _GEN_2390; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2586 = _T_23 ? plru2_16 : _GEN_2391; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2587 = _T_23 ? plru2_17 : _GEN_2392; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2588 = _T_23 ? plru2_18 : _GEN_2393; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2589 = _T_23 ? plru2_19 : _GEN_2394; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2590 = _T_23 ? plru2_20 : _GEN_2395; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2591 = _T_23 ? plru2_21 : _GEN_2396; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2592 = _T_23 ? plru2_22 : _GEN_2397; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2593 = _T_23 ? plru2_23 : _GEN_2398; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2594 = _T_23 ? plru2_24 : _GEN_2399; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2595 = _T_23 ? plru2_25 : _GEN_2400; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2596 = _T_23 ? plru2_26 : _GEN_2401; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2597 = _T_23 ? plru2_27 : _GEN_2402; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2598 = _T_23 ? plru2_28 : _GEN_2403; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2599 = _T_23 ? plru2_29 : _GEN_2404; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2600 = _T_23 ? plru2_30 : _GEN_2405; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2601 = _T_23 ? plru2_31 : _GEN_2406; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2602 = _T_23 ? plru2_32 : _GEN_2407; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2603 = _T_23 ? plru2_33 : _GEN_2408; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2604 = _T_23 ? plru2_34 : _GEN_2409; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2605 = _T_23 ? plru2_35 : _GEN_2410; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2606 = _T_23 ? plru2_36 : _GEN_2411; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2607 = _T_23 ? plru2_37 : _GEN_2412; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2608 = _T_23 ? plru2_38 : _GEN_2413; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2609 = _T_23 ? plru2_39 : _GEN_2414; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2610 = _T_23 ? plru2_40 : _GEN_2415; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2611 = _T_23 ? plru2_41 : _GEN_2416; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2612 = _T_23 ? plru2_42 : _GEN_2417; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2613 = _T_23 ? plru2_43 : _GEN_2418; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2614 = _T_23 ? plru2_44 : _GEN_2419; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2615 = _T_23 ? plru2_45 : _GEN_2420; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2616 = _T_23 ? plru2_46 : _GEN_2421; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2617 = _T_23 ? plru2_47 : _GEN_2422; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2618 = _T_23 ? plru2_48 : _GEN_2423; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2619 = _T_23 ? plru2_49 : _GEN_2424; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2620 = _T_23 ? plru2_50 : _GEN_2425; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2621 = _T_23 ? plru2_51 : _GEN_2426; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2622 = _T_23 ? plru2_52 : _GEN_2427; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2623 = _T_23 ? plru2_53 : _GEN_2428; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2624 = _T_23 ? plru2_54 : _GEN_2429; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2625 = _T_23 ? plru2_55 : _GEN_2430; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2626 = _T_23 ? plru2_56 : _GEN_2431; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2627 = _T_23 ? plru2_57 : _GEN_2432; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2628 = _T_23 ? plru2_58 : _GEN_2433; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2629 = _T_23 ? plru2_59 : _GEN_2434; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2630 = _T_23 ? plru2_60 : _GEN_2435; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2631 = _T_23 ? plru2_61 : _GEN_2436; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2632 = _T_23 ? plru2_62 : _GEN_2437; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire  _GEN_2633 = _T_23 ? plru2_63 : _GEN_2438; // @[Conditional.scala 39:67 Cache.scala 135:22]
  wire [63:0] _GEN_2634 = _T_23 ? 64'h0 : _GEN_2439; // @[Conditional.scala 39:67 Cache.scala 277:22]
  wire  _GEN_2635 = _T_16 ? _GEN_992 : fi_ready; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2637 = _T_16 ? _GEN_994 : _GEN_3; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2638 = _T_16 ? _GEN_995 : 128'h0; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_2639 = _T_16 ? _GEN_996 : 21'h0; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_2641 = _T_16 ? _GEN_999 : fi_ready; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2643 = _T_16 ? _GEN_1001 : _GEN_3; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2644 = _T_16 ? _GEN_1002 : 128'h0; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_2645 = _T_16 ? _GEN_1003 : 21'h0; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_2647 = _T_16 ? _GEN_1006 : fi_ready; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2649 = _T_16 ? _GEN_1008 : _GEN_3; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2650 = _T_16 ? _GEN_1009 : 128'h0; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_2651 = _T_16 ? _GEN_1010 : 21'h0; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_2653 = _T_16 ? _GEN_1013 : fi_ready; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2655 = _T_16 ? _GEN_1015 : _GEN_3; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2656 = _T_16 ? _GEN_1016 : 128'h0; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_2657 = _T_16 ? _GEN_1017 : 21'h0; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire [3:0] _GEN_2659 = _T_16 ? _GEN_1339 : _GEN_2440; // @[Conditional.scala 39:67]
  wire  _GEN_2660 = _T_16 ? _GEN_1340 : _GEN_2442; // @[Conditional.scala 39:67]
  wire  _GEN_2661 = _T_16 ? _GEN_1341 : _GEN_2443; // @[Conditional.scala 39:67]
  wire  _GEN_2662 = _T_16 ? _GEN_1342 : _GEN_2444; // @[Conditional.scala 39:67]
  wire  _GEN_2663 = _T_16 ? _GEN_1343 : _GEN_2445; // @[Conditional.scala 39:67]
  wire  _GEN_2664 = _T_16 ? _GEN_1344 : _GEN_2446; // @[Conditional.scala 39:67]
  wire  _GEN_2665 = _T_16 ? _GEN_1345 : _GEN_2447; // @[Conditional.scala 39:67]
  wire  _GEN_2666 = _T_16 ? _GEN_1346 : _GEN_2448; // @[Conditional.scala 39:67]
  wire  _GEN_2667 = _T_16 ? _GEN_1347 : _GEN_2449; // @[Conditional.scala 39:67]
  wire  _GEN_2668 = _T_16 ? _GEN_1348 : _GEN_2450; // @[Conditional.scala 39:67]
  wire  _GEN_2669 = _T_16 ? _GEN_1349 : _GEN_2451; // @[Conditional.scala 39:67]
  wire  _GEN_2670 = _T_16 ? _GEN_1350 : _GEN_2452; // @[Conditional.scala 39:67]
  wire  _GEN_2671 = _T_16 ? _GEN_1351 : _GEN_2453; // @[Conditional.scala 39:67]
  wire  _GEN_2672 = _T_16 ? _GEN_1352 : _GEN_2454; // @[Conditional.scala 39:67]
  wire  _GEN_2673 = _T_16 ? _GEN_1353 : _GEN_2455; // @[Conditional.scala 39:67]
  wire  _GEN_2674 = _T_16 ? _GEN_1354 : _GEN_2456; // @[Conditional.scala 39:67]
  wire  _GEN_2675 = _T_16 ? _GEN_1355 : _GEN_2457; // @[Conditional.scala 39:67]
  wire  _GEN_2676 = _T_16 ? _GEN_1356 : _GEN_2458; // @[Conditional.scala 39:67]
  wire  _GEN_2677 = _T_16 ? _GEN_1357 : _GEN_2459; // @[Conditional.scala 39:67]
  wire  _GEN_2678 = _T_16 ? _GEN_1358 : _GEN_2460; // @[Conditional.scala 39:67]
  wire  _GEN_2679 = _T_16 ? _GEN_1359 : _GEN_2461; // @[Conditional.scala 39:67]
  wire  _GEN_2680 = _T_16 ? _GEN_1360 : _GEN_2462; // @[Conditional.scala 39:67]
  wire  _GEN_2681 = _T_16 ? _GEN_1361 : _GEN_2463; // @[Conditional.scala 39:67]
  wire  _GEN_2682 = _T_16 ? _GEN_1362 : _GEN_2464; // @[Conditional.scala 39:67]
  wire  _GEN_2683 = _T_16 ? _GEN_1363 : _GEN_2465; // @[Conditional.scala 39:67]
  wire  _GEN_2684 = _T_16 ? _GEN_1364 : _GEN_2466; // @[Conditional.scala 39:67]
  wire  _GEN_2685 = _T_16 ? _GEN_1365 : _GEN_2467; // @[Conditional.scala 39:67]
  wire  _GEN_2686 = _T_16 ? _GEN_1366 : _GEN_2468; // @[Conditional.scala 39:67]
  wire  _GEN_2687 = _T_16 ? _GEN_1367 : _GEN_2469; // @[Conditional.scala 39:67]
  wire  _GEN_2688 = _T_16 ? _GEN_1368 : _GEN_2470; // @[Conditional.scala 39:67]
  wire  _GEN_2689 = _T_16 ? _GEN_1369 : _GEN_2471; // @[Conditional.scala 39:67]
  wire  _GEN_2690 = _T_16 ? _GEN_1370 : _GEN_2472; // @[Conditional.scala 39:67]
  wire  _GEN_2691 = _T_16 ? _GEN_1371 : _GEN_2473; // @[Conditional.scala 39:67]
  wire  _GEN_2692 = _T_16 ? _GEN_1372 : _GEN_2474; // @[Conditional.scala 39:67]
  wire  _GEN_2693 = _T_16 ? _GEN_1373 : _GEN_2475; // @[Conditional.scala 39:67]
  wire  _GEN_2694 = _T_16 ? _GEN_1374 : _GEN_2476; // @[Conditional.scala 39:67]
  wire  _GEN_2695 = _T_16 ? _GEN_1375 : _GEN_2477; // @[Conditional.scala 39:67]
  wire  _GEN_2696 = _T_16 ? _GEN_1376 : _GEN_2478; // @[Conditional.scala 39:67]
  wire  _GEN_2697 = _T_16 ? _GEN_1377 : _GEN_2479; // @[Conditional.scala 39:67]
  wire  _GEN_2698 = _T_16 ? _GEN_1378 : _GEN_2480; // @[Conditional.scala 39:67]
  wire  _GEN_2699 = _T_16 ? _GEN_1379 : _GEN_2481; // @[Conditional.scala 39:67]
  wire  _GEN_2700 = _T_16 ? _GEN_1380 : _GEN_2482; // @[Conditional.scala 39:67]
  wire  _GEN_2701 = _T_16 ? _GEN_1381 : _GEN_2483; // @[Conditional.scala 39:67]
  wire  _GEN_2702 = _T_16 ? _GEN_1382 : _GEN_2484; // @[Conditional.scala 39:67]
  wire  _GEN_2703 = _T_16 ? _GEN_1383 : _GEN_2485; // @[Conditional.scala 39:67]
  wire  _GEN_2704 = _T_16 ? _GEN_1384 : _GEN_2486; // @[Conditional.scala 39:67]
  wire  _GEN_2705 = _T_16 ? _GEN_1385 : _GEN_2487; // @[Conditional.scala 39:67]
  wire  _GEN_2706 = _T_16 ? _GEN_1386 : _GEN_2488; // @[Conditional.scala 39:67]
  wire  _GEN_2707 = _T_16 ? _GEN_1387 : _GEN_2489; // @[Conditional.scala 39:67]
  wire  _GEN_2708 = _T_16 ? _GEN_1388 : _GEN_2490; // @[Conditional.scala 39:67]
  wire  _GEN_2709 = _T_16 ? _GEN_1389 : _GEN_2491; // @[Conditional.scala 39:67]
  wire  _GEN_2710 = _T_16 ? _GEN_1390 : _GEN_2492; // @[Conditional.scala 39:67]
  wire  _GEN_2711 = _T_16 ? _GEN_1391 : _GEN_2493; // @[Conditional.scala 39:67]
  wire  _GEN_2712 = _T_16 ? _GEN_1392 : _GEN_2494; // @[Conditional.scala 39:67]
  wire  _GEN_2713 = _T_16 ? _GEN_1393 : _GEN_2495; // @[Conditional.scala 39:67]
  wire  _GEN_2714 = _T_16 ? _GEN_1394 : _GEN_2496; // @[Conditional.scala 39:67]
  wire  _GEN_2715 = _T_16 ? _GEN_1395 : _GEN_2497; // @[Conditional.scala 39:67]
  wire  _GEN_2716 = _T_16 ? _GEN_1396 : _GEN_2498; // @[Conditional.scala 39:67]
  wire  _GEN_2717 = _T_16 ? _GEN_1397 : _GEN_2499; // @[Conditional.scala 39:67]
  wire  _GEN_2718 = _T_16 ? _GEN_1398 : _GEN_2500; // @[Conditional.scala 39:67]
  wire  _GEN_2719 = _T_16 ? _GEN_1399 : _GEN_2501; // @[Conditional.scala 39:67]
  wire  _GEN_2720 = _T_16 ? _GEN_1400 : _GEN_2502; // @[Conditional.scala 39:67]
  wire  _GEN_2721 = _T_16 ? _GEN_1401 : _GEN_2503; // @[Conditional.scala 39:67]
  wire  _GEN_2722 = _T_16 ? _GEN_1402 : _GEN_2504; // @[Conditional.scala 39:67]
  wire  _GEN_2723 = _T_16 ? _GEN_1403 : _GEN_2505; // @[Conditional.scala 39:67]
  wire  _GEN_2724 = _T_16 ? _GEN_1404 : _GEN_2506; // @[Conditional.scala 39:67]
  wire  _GEN_2725 = _T_16 ? _GEN_1405 : _GEN_2507; // @[Conditional.scala 39:67]
  wire  _GEN_2726 = _T_16 ? _GEN_1406 : _GEN_2508; // @[Conditional.scala 39:67]
  wire  _GEN_2727 = _T_16 ? _GEN_1407 : _GEN_2509; // @[Conditional.scala 39:67]
  wire  _GEN_2728 = _T_16 ? _GEN_1408 : _GEN_2510; // @[Conditional.scala 39:67]
  wire  _GEN_2729 = _T_16 ? _GEN_1409 : _GEN_2511; // @[Conditional.scala 39:67]
  wire  _GEN_2730 = _T_16 ? _GEN_1410 : _GEN_2512; // @[Conditional.scala 39:67]
  wire  _GEN_2731 = _T_16 ? _GEN_1411 : _GEN_2513; // @[Conditional.scala 39:67]
  wire  _GEN_2732 = _T_16 ? _GEN_1412 : _GEN_2514; // @[Conditional.scala 39:67]
  wire  _GEN_2733 = _T_16 ? _GEN_1413 : _GEN_2515; // @[Conditional.scala 39:67]
  wire  _GEN_2734 = _T_16 ? _GEN_1414 : _GEN_2516; // @[Conditional.scala 39:67]
  wire  _GEN_2735 = _T_16 ? _GEN_1415 : _GEN_2517; // @[Conditional.scala 39:67]
  wire  _GEN_2736 = _T_16 ? _GEN_1416 : _GEN_2518; // @[Conditional.scala 39:67]
  wire  _GEN_2737 = _T_16 ? _GEN_1417 : _GEN_2519; // @[Conditional.scala 39:67]
  wire  _GEN_2738 = _T_16 ? _GEN_1418 : _GEN_2520; // @[Conditional.scala 39:67]
  wire  _GEN_2739 = _T_16 ? _GEN_1419 : _GEN_2521; // @[Conditional.scala 39:67]
  wire  _GEN_2740 = _T_16 ? _GEN_1420 : _GEN_2522; // @[Conditional.scala 39:67]
  wire  _GEN_2741 = _T_16 ? _GEN_1421 : _GEN_2523; // @[Conditional.scala 39:67]
  wire  _GEN_2742 = _T_16 ? _GEN_1422 : _GEN_2524; // @[Conditional.scala 39:67]
  wire  _GEN_2743 = _T_16 ? _GEN_1423 : _GEN_2525; // @[Conditional.scala 39:67]
  wire  _GEN_2744 = _T_16 ? _GEN_1424 : _GEN_2526; // @[Conditional.scala 39:67]
  wire  _GEN_2745 = _T_16 ? _GEN_1425 : _GEN_2527; // @[Conditional.scala 39:67]
  wire  _GEN_2746 = _T_16 ? _GEN_1426 : _GEN_2528; // @[Conditional.scala 39:67]
  wire  _GEN_2747 = _T_16 ? _GEN_1427 : _GEN_2529; // @[Conditional.scala 39:67]
  wire  _GEN_2748 = _T_16 ? _GEN_1428 : _GEN_2530; // @[Conditional.scala 39:67]
  wire  _GEN_2749 = _T_16 ? _GEN_1429 : _GEN_2531; // @[Conditional.scala 39:67]
  wire  _GEN_2750 = _T_16 ? _GEN_1430 : _GEN_2532; // @[Conditional.scala 39:67]
  wire  _GEN_2751 = _T_16 ? _GEN_1431 : _GEN_2533; // @[Conditional.scala 39:67]
  wire  _GEN_2752 = _T_16 ? _GEN_1432 : _GEN_2534; // @[Conditional.scala 39:67]
  wire  _GEN_2753 = _T_16 ? _GEN_1433 : _GEN_2535; // @[Conditional.scala 39:67]
  wire  _GEN_2754 = _T_16 ? _GEN_1434 : _GEN_2536; // @[Conditional.scala 39:67]
  wire  _GEN_2755 = _T_16 ? _GEN_1435 : _GEN_2537; // @[Conditional.scala 39:67]
  wire  _GEN_2756 = _T_16 ? _GEN_1436 : _GEN_2538; // @[Conditional.scala 39:67]
  wire  _GEN_2757 = _T_16 ? _GEN_1437 : _GEN_2539; // @[Conditional.scala 39:67]
  wire  _GEN_2758 = _T_16 ? _GEN_1438 : _GEN_2540; // @[Conditional.scala 39:67]
  wire  _GEN_2759 = _T_16 ? _GEN_1439 : _GEN_2541; // @[Conditional.scala 39:67]
  wire  _GEN_2760 = _T_16 ? _GEN_1440 : _GEN_2542; // @[Conditional.scala 39:67]
  wire  _GEN_2761 = _T_16 ? _GEN_1441 : _GEN_2543; // @[Conditional.scala 39:67]
  wire  _GEN_2762 = _T_16 ? _GEN_1442 : _GEN_2544; // @[Conditional.scala 39:67]
  wire  _GEN_2763 = _T_16 ? _GEN_1443 : _GEN_2545; // @[Conditional.scala 39:67]
  wire  _GEN_2764 = _T_16 ? _GEN_1444 : _GEN_2546; // @[Conditional.scala 39:67]
  wire  _GEN_2765 = _T_16 ? _GEN_1445 : _GEN_2547; // @[Conditional.scala 39:67]
  wire  _GEN_2766 = _T_16 ? _GEN_1446 : _GEN_2548; // @[Conditional.scala 39:67]
  wire  _GEN_2767 = _T_16 ? _GEN_1447 : _GEN_2549; // @[Conditional.scala 39:67]
  wire  _GEN_2768 = _T_16 ? _GEN_1448 : _GEN_2550; // @[Conditional.scala 39:67]
  wire  _GEN_2769 = _T_16 ? _GEN_1449 : _GEN_2551; // @[Conditional.scala 39:67]
  wire  _GEN_2770 = _T_16 ? _GEN_1450 : _GEN_2552; // @[Conditional.scala 39:67]
  wire  _GEN_2771 = _T_16 ? _GEN_1451 : _GEN_2553; // @[Conditional.scala 39:67]
  wire  _GEN_2772 = _T_16 ? _GEN_1452 : _GEN_2554; // @[Conditional.scala 39:67]
  wire  _GEN_2773 = _T_16 ? _GEN_1453 : _GEN_2555; // @[Conditional.scala 39:67]
  wire  _GEN_2774 = _T_16 ? _GEN_1454 : _GEN_2556; // @[Conditional.scala 39:67]
  wire  _GEN_2775 = _T_16 ? _GEN_1455 : _GEN_2557; // @[Conditional.scala 39:67]
  wire  _GEN_2776 = _T_16 ? _GEN_1456 : _GEN_2558; // @[Conditional.scala 39:67]
  wire  _GEN_2777 = _T_16 ? _GEN_1457 : _GEN_2559; // @[Conditional.scala 39:67]
  wire  _GEN_2778 = _T_16 ? _GEN_1458 : _GEN_2560; // @[Conditional.scala 39:67]
  wire  _GEN_2779 = _T_16 ? _GEN_1459 : _GEN_2561; // @[Conditional.scala 39:67]
  wire  _GEN_2780 = _T_16 ? _GEN_1460 : _GEN_2562; // @[Conditional.scala 39:67]
  wire  _GEN_2781 = _T_16 ? _GEN_1461 : _GEN_2563; // @[Conditional.scala 39:67]
  wire  _GEN_2782 = _T_16 ? _GEN_1462 : _GEN_2564; // @[Conditional.scala 39:67]
  wire  _GEN_2783 = _T_16 ? _GEN_1463 : _GEN_2565; // @[Conditional.scala 39:67]
  wire  _GEN_2784 = _T_16 ? _GEN_1464 : _GEN_2566; // @[Conditional.scala 39:67]
  wire  _GEN_2785 = _T_16 ? _GEN_1465 : _GEN_2567; // @[Conditional.scala 39:67]
  wire  _GEN_2786 = _T_16 ? _GEN_1466 : _GEN_2568; // @[Conditional.scala 39:67]
  wire  _GEN_2787 = _T_16 ? _GEN_1467 : _GEN_2569; // @[Conditional.scala 39:67]
  wire  _GEN_2788 = _T_16 ? _GEN_1468 : _GEN_2570; // @[Conditional.scala 39:67]
  wire  _GEN_2789 = _T_16 ? _GEN_1469 : _GEN_2571; // @[Conditional.scala 39:67]
  wire  _GEN_2790 = _T_16 ? _GEN_1470 : _GEN_2572; // @[Conditional.scala 39:67]
  wire  _GEN_2791 = _T_16 ? _GEN_1471 : _GEN_2573; // @[Conditional.scala 39:67]
  wire  _GEN_2792 = _T_16 ? _GEN_1472 : _GEN_2574; // @[Conditional.scala 39:67]
  wire  _GEN_2793 = _T_16 ? _GEN_1473 : _GEN_2575; // @[Conditional.scala 39:67]
  wire  _GEN_2794 = _T_16 ? _GEN_1474 : _GEN_2576; // @[Conditional.scala 39:67]
  wire  _GEN_2795 = _T_16 ? _GEN_1475 : _GEN_2577; // @[Conditional.scala 39:67]
  wire  _GEN_2796 = _T_16 ? _GEN_1476 : _GEN_2578; // @[Conditional.scala 39:67]
  wire  _GEN_2797 = _T_16 ? _GEN_1477 : _GEN_2579; // @[Conditional.scala 39:67]
  wire  _GEN_2798 = _T_16 ? _GEN_1478 : _GEN_2580; // @[Conditional.scala 39:67]
  wire  _GEN_2799 = _T_16 ? _GEN_1479 : _GEN_2581; // @[Conditional.scala 39:67]
  wire  _GEN_2800 = _T_16 ? _GEN_1480 : _GEN_2582; // @[Conditional.scala 39:67]
  wire  _GEN_2801 = _T_16 ? _GEN_1481 : _GEN_2583; // @[Conditional.scala 39:67]
  wire  _GEN_2802 = _T_16 ? _GEN_1482 : _GEN_2584; // @[Conditional.scala 39:67]
  wire  _GEN_2803 = _T_16 ? _GEN_1483 : _GEN_2585; // @[Conditional.scala 39:67]
  wire  _GEN_2804 = _T_16 ? _GEN_1484 : _GEN_2586; // @[Conditional.scala 39:67]
  wire  _GEN_2805 = _T_16 ? _GEN_1485 : _GEN_2587; // @[Conditional.scala 39:67]
  wire  _GEN_2806 = _T_16 ? _GEN_1486 : _GEN_2588; // @[Conditional.scala 39:67]
  wire  _GEN_2807 = _T_16 ? _GEN_1487 : _GEN_2589; // @[Conditional.scala 39:67]
  wire  _GEN_2808 = _T_16 ? _GEN_1488 : _GEN_2590; // @[Conditional.scala 39:67]
  wire  _GEN_2809 = _T_16 ? _GEN_1489 : _GEN_2591; // @[Conditional.scala 39:67]
  wire  _GEN_2810 = _T_16 ? _GEN_1490 : _GEN_2592; // @[Conditional.scala 39:67]
  wire  _GEN_2811 = _T_16 ? _GEN_1491 : _GEN_2593; // @[Conditional.scala 39:67]
  wire  _GEN_2812 = _T_16 ? _GEN_1492 : _GEN_2594; // @[Conditional.scala 39:67]
  wire  _GEN_2813 = _T_16 ? _GEN_1493 : _GEN_2595; // @[Conditional.scala 39:67]
  wire  _GEN_2814 = _T_16 ? _GEN_1494 : _GEN_2596; // @[Conditional.scala 39:67]
  wire  _GEN_2815 = _T_16 ? _GEN_1495 : _GEN_2597; // @[Conditional.scala 39:67]
  wire  _GEN_2816 = _T_16 ? _GEN_1496 : _GEN_2598; // @[Conditional.scala 39:67]
  wire  _GEN_2817 = _T_16 ? _GEN_1497 : _GEN_2599; // @[Conditional.scala 39:67]
  wire  _GEN_2818 = _T_16 ? _GEN_1498 : _GEN_2600; // @[Conditional.scala 39:67]
  wire  _GEN_2819 = _T_16 ? _GEN_1499 : _GEN_2601; // @[Conditional.scala 39:67]
  wire  _GEN_2820 = _T_16 ? _GEN_1500 : _GEN_2602; // @[Conditional.scala 39:67]
  wire  _GEN_2821 = _T_16 ? _GEN_1501 : _GEN_2603; // @[Conditional.scala 39:67]
  wire  _GEN_2822 = _T_16 ? _GEN_1502 : _GEN_2604; // @[Conditional.scala 39:67]
  wire  _GEN_2823 = _T_16 ? _GEN_1503 : _GEN_2605; // @[Conditional.scala 39:67]
  wire  _GEN_2824 = _T_16 ? _GEN_1504 : _GEN_2606; // @[Conditional.scala 39:67]
  wire  _GEN_2825 = _T_16 ? _GEN_1505 : _GEN_2607; // @[Conditional.scala 39:67]
  wire  _GEN_2826 = _T_16 ? _GEN_1506 : _GEN_2608; // @[Conditional.scala 39:67]
  wire  _GEN_2827 = _T_16 ? _GEN_1507 : _GEN_2609; // @[Conditional.scala 39:67]
  wire  _GEN_2828 = _T_16 ? _GEN_1508 : _GEN_2610; // @[Conditional.scala 39:67]
  wire  _GEN_2829 = _T_16 ? _GEN_1509 : _GEN_2611; // @[Conditional.scala 39:67]
  wire  _GEN_2830 = _T_16 ? _GEN_1510 : _GEN_2612; // @[Conditional.scala 39:67]
  wire  _GEN_2831 = _T_16 ? _GEN_1511 : _GEN_2613; // @[Conditional.scala 39:67]
  wire  _GEN_2832 = _T_16 ? _GEN_1512 : _GEN_2614; // @[Conditional.scala 39:67]
  wire  _GEN_2833 = _T_16 ? _GEN_1513 : _GEN_2615; // @[Conditional.scala 39:67]
  wire  _GEN_2834 = _T_16 ? _GEN_1514 : _GEN_2616; // @[Conditional.scala 39:67]
  wire  _GEN_2835 = _T_16 ? _GEN_1515 : _GEN_2617; // @[Conditional.scala 39:67]
  wire  _GEN_2836 = _T_16 ? _GEN_1516 : _GEN_2618; // @[Conditional.scala 39:67]
  wire  _GEN_2837 = _T_16 ? _GEN_1517 : _GEN_2619; // @[Conditional.scala 39:67]
  wire  _GEN_2838 = _T_16 ? _GEN_1518 : _GEN_2620; // @[Conditional.scala 39:67]
  wire  _GEN_2839 = _T_16 ? _GEN_1519 : _GEN_2621; // @[Conditional.scala 39:67]
  wire  _GEN_2840 = _T_16 ? _GEN_1520 : _GEN_2622; // @[Conditional.scala 39:67]
  wire  _GEN_2841 = _T_16 ? _GEN_1521 : _GEN_2623; // @[Conditional.scala 39:67]
  wire  _GEN_2842 = _T_16 ? _GEN_1522 : _GEN_2624; // @[Conditional.scala 39:67]
  wire  _GEN_2843 = _T_16 ? _GEN_1523 : _GEN_2625; // @[Conditional.scala 39:67]
  wire  _GEN_2844 = _T_16 ? _GEN_1524 : _GEN_2626; // @[Conditional.scala 39:67]
  wire  _GEN_2845 = _T_16 ? _GEN_1525 : _GEN_2627; // @[Conditional.scala 39:67]
  wire  _GEN_2846 = _T_16 ? _GEN_1526 : _GEN_2628; // @[Conditional.scala 39:67]
  wire  _GEN_2847 = _T_16 ? _GEN_1527 : _GEN_2629; // @[Conditional.scala 39:67]
  wire  _GEN_2848 = _T_16 ? _GEN_1528 : _GEN_2630; // @[Conditional.scala 39:67]
  wire  _GEN_2849 = _T_16 ? _GEN_1529 : _GEN_2631; // @[Conditional.scala 39:67]
  wire  _GEN_2850 = _T_16 ? _GEN_1530 : _GEN_2632; // @[Conditional.scala 39:67]
  wire  _GEN_2851 = _T_16 ? _GEN_1531 : _GEN_2633; // @[Conditional.scala 39:67]
  wire  _GEN_2852 = _T_16 ? _GEN_27 : _GEN_2441; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_2853 = _T_16 ? 64'h0 : _GEN_2634; // @[Conditional.scala 39:67 Cache.scala 277:22]
  wire [3:0] _GEN_2856 = _T_13 ? _GEN_990 : _GEN_2659; // @[Conditional.scala 39:67]
  wire  _GEN_2857 = _T_13 ? fi_ready : _GEN_2635; // @[Conditional.scala 39:67]
  wire  _GEN_2858 = _T_13 ? 1'h0 : _T_16 & _T_17; // @[Conditional.scala 39:67 Cache.scala 110:14]
  wire [5:0] _GEN_2859 = _T_13 ? _GEN_3 : _GEN_2637; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2860 = _T_13 ? 128'h0 : _GEN_2638; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_2861 = _T_13 ? 21'h0 : _GEN_2639; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_2862 = _T_13 ? 1'h0 : _T_16 & _GEN_997; // @[Conditional.scala 39:67 Cache.scala 118:18]
  wire  _GEN_2863 = _T_13 ? fi_ready : _GEN_2641; // @[Conditional.scala 39:67]
  wire  _GEN_2864 = _T_13 ? 1'h0 : _T_16 & _T_18; // @[Conditional.scala 39:67 Cache.scala 110:14]
  wire [5:0] _GEN_2865 = _T_13 ? _GEN_3 : _GEN_2643; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2866 = _T_13 ? 128'h0 : _GEN_2644; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_2867 = _T_13 ? 21'h0 : _GEN_2645; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_2868 = _T_13 ? 1'h0 : _T_16 & _GEN_1004; // @[Conditional.scala 39:67 Cache.scala 118:18]
  wire  _GEN_2869 = _T_13 ? fi_ready : _GEN_2647; // @[Conditional.scala 39:67]
  wire  _GEN_2870 = _T_13 ? 1'h0 : _T_16 & _T_19; // @[Conditional.scala 39:67 Cache.scala 110:14]
  wire [5:0] _GEN_2871 = _T_13 ? _GEN_3 : _GEN_2649; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2872 = _T_13 ? 128'h0 : _GEN_2650; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_2873 = _T_13 ? 21'h0 : _GEN_2651; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_2874 = _T_13 ? 1'h0 : _T_16 & _GEN_1011; // @[Conditional.scala 39:67 Cache.scala 118:18]
  wire  _GEN_2875 = _T_13 ? fi_ready : _GEN_2653; // @[Conditional.scala 39:67]
  wire  _GEN_2876 = _T_13 ? 1'h0 : _T_16 & _T_20; // @[Conditional.scala 39:67 Cache.scala 110:14]
  wire [5:0] _GEN_2877 = _T_13 ? _GEN_3 : _GEN_2655; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2878 = _T_13 ? 128'h0 : _GEN_2656; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_2879 = _T_13 ? 21'h0 : _GEN_2657; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_2880 = _T_13 ? 1'h0 : _T_16 & _GEN_1018; // @[Conditional.scala 39:67 Cache.scala 118:18]
  wire [63:0] _GEN_3074 = _T_13 ? 64'h0 : _GEN_2853; // @[Conditional.scala 39:67 Cache.scala 277:22]
  wire [3:0] _GEN_3075 = _T_11 ? _GEN_984 : _GEN_2856; // @[Conditional.scala 39:67]
  wire  _GEN_3078 = _T_11 ? fi_ready : _GEN_2857; // @[Conditional.scala 39:67]
  wire  _GEN_3079 = _T_11 ? 1'h0 : _GEN_2858; // @[Conditional.scala 39:67 Cache.scala 110:14]
  wire [5:0] _GEN_3080 = _T_11 ? _GEN_3 : _GEN_2859; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_3081 = _T_11 ? 128'h0 : _GEN_2860; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_3082 = _T_11 ? 21'h0 : _GEN_2861; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_3083 = _T_11 ? 1'h0 : _GEN_2862; // @[Conditional.scala 39:67 Cache.scala 118:18]
  wire  _GEN_3084 = _T_11 ? fi_ready : _GEN_2863; // @[Conditional.scala 39:67]
  wire  _GEN_3085 = _T_11 ? 1'h0 : _GEN_2864; // @[Conditional.scala 39:67 Cache.scala 110:14]
  wire [5:0] _GEN_3086 = _T_11 ? _GEN_3 : _GEN_2865; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_3087 = _T_11 ? 128'h0 : _GEN_2866; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_3088 = _T_11 ? 21'h0 : _GEN_2867; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_3089 = _T_11 ? 1'h0 : _GEN_2868; // @[Conditional.scala 39:67 Cache.scala 118:18]
  wire  _GEN_3090 = _T_11 ? fi_ready : _GEN_2869; // @[Conditional.scala 39:67]
  wire  _GEN_3091 = _T_11 ? 1'h0 : _GEN_2870; // @[Conditional.scala 39:67 Cache.scala 110:14]
  wire [5:0] _GEN_3092 = _T_11 ? _GEN_3 : _GEN_2871; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_3093 = _T_11 ? 128'h0 : _GEN_2872; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_3094 = _T_11 ? 21'h0 : _GEN_2873; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_3095 = _T_11 ? 1'h0 : _GEN_2874; // @[Conditional.scala 39:67 Cache.scala 118:18]
  wire  _GEN_3096 = _T_11 ? fi_ready : _GEN_2875; // @[Conditional.scala 39:67]
  wire  _GEN_3097 = _T_11 ? 1'h0 : _GEN_2876; // @[Conditional.scala 39:67 Cache.scala 110:14]
  wire [5:0] _GEN_3098 = _T_11 ? _GEN_3 : _GEN_2877; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_3099 = _T_11 ? 128'h0 : _GEN_2878; // @[Conditional.scala 39:67 Cache.scala 112:16]
  wire [20:0] _GEN_3100 = _T_11 ? 21'h0 : _GEN_2879; // @[Conditional.scala 39:67 Cache.scala 116:16]
  wire  _GEN_3101 = _T_11 ? 1'h0 : _GEN_2880; // @[Conditional.scala 39:67 Cache.scala 118:18]
  wire [63:0] _GEN_3295 = _T_11 ? 64'h0 : _GEN_3074; // @[Conditional.scala 39:67 Cache.scala 277:22]
  wire  _GEN_3489 = _T_2 ? _GEN_967 : _GEN_3078; // @[Conditional.scala 40:58]
  wire [5:0] _GEN_3491 = _T_2 ? _GEN_969 : _GEN_3080; // @[Conditional.scala 40:58]
  wire  _GEN_3494 = _T_2 ? _GEN_971 : _GEN_3084; // @[Conditional.scala 40:58]
  wire [5:0] _GEN_3496 = _T_2 ? _GEN_973 : _GEN_3086; // @[Conditional.scala 40:58]
  wire  _GEN_3499 = _T_2 ? _GEN_975 : _GEN_3090; // @[Conditional.scala 40:58]
  wire [5:0] _GEN_3501 = _T_2 ? _GEN_977 : _GEN_3092; // @[Conditional.scala 40:58]
  wire  _GEN_3504 = _T_2 ? _GEN_979 : _GEN_3096; // @[Conditional.scala 40:58]
  wire [5:0] _GEN_3506 = _T_2 ? _GEN_981 : _GEN_3098; // @[Conditional.scala 40:58]
  reg [7:0] fi_counter; // @[Cache.scala 402:27]
  wire [1:0] fi_sram_idx = fi_counter[7:6]; // @[Cache.scala 403:31]
  wire [5:0] fi_line_idx = fi_counter[5:0]; // @[Cache.scala 404:31]
  wire  _fi_update_T = fi_state == 3'h2; // @[Cache.scala 407:29]
  wire  _fi_update_T_1 = fi_state == 3'h1; // @[Cache.scala 407:65]
  reg  fi_update_REG; // @[Cache.scala 407:55]
  wire  fi_update = fi_state == 3'h2 & fi_update_REG; // @[Cache.scala 407:44]
  reg [127:0] fi_wdata_r; // @[Reg.scala 27:20]
  wire [127:0] _GEN_3523 = 2'h1 == fi_sram_idx ? sram_out_1 : sram_out_0; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [127:0] _GEN_3524 = 2'h2 == fi_sram_idx ? sram_out_2 : _GEN_3523; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [127:0] _GEN_3525 = 2'h3 == fi_sram_idx ? sram_out_3 : _GEN_3524; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [127:0] _GEN_3526 = fi_update ? _GEN_3525 : fi_wdata_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  reg [20:0] fi_tag_r; // @[Reg.scala 27:20]
  wire [20:0] _GEN_3528 = 2'h1 == fi_sram_idx ? tag_out_1 : tag_out_0; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [20:0] _GEN_3529 = 2'h2 == fi_sram_idx ? tag_out_2 : _GEN_3528; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [20:0] _GEN_3530 = 2'h3 == fi_sram_idx ? tag_out_3 : _GEN_3529; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [20:0] _GEN_3531 = fi_update ? _GEN_3530 : fi_tag_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [7:0] fi_counter_next = fi_counter + 8'h1; // @[Cache.scala 435:38]
  wire [5:0] _GEN_3534 = _fi_update_T_1 ? fi_line_idx : _GEN_3491; // @[Cache.scala 437:40 Cache.scala 440:19]
  wire [5:0] _GEN_3536 = _fi_update_T_1 ? fi_line_idx : _GEN_3496; // @[Cache.scala 437:40 Cache.scala 440:19]
  wire [5:0] _GEN_3538 = _fi_update_T_1 ? fi_line_idx : _GEN_3501; // @[Cache.scala 437:40 Cache.scala 440:19]
  wire [5:0] _GEN_3540 = _fi_update_T_1 ? fi_line_idx : _GEN_3506; // @[Cache.scala 437:40 Cache.scala 440:19]
  wire [5:0] _GEN_3543 = fi_sram_idx == 2'h0 ? fi_line_idx : _GEN_3534; // @[Cache.scala 457:38 Cache.scala 458:28]
  wire [5:0] _GEN_3545 = fi_sram_idx == 2'h1 ? fi_line_idx : _GEN_3536; // @[Cache.scala 457:38 Cache.scala 458:28]
  wire  _GEN_3546 = fi_sram_idx == 2'h1 ? meta_1_io_valid_r_async & meta_1_io_dirty_r_async : fi_sram_idx == 2'h0 & (
    meta_0_io_valid_r_async & meta_0_io_dirty_r_async); // @[Cache.scala 457:38 Cache.scala 459:22]
  wire [5:0] _GEN_3547 = fi_sram_idx == 2'h2 ? fi_line_idx : _GEN_3538; // @[Cache.scala 457:38 Cache.scala 458:28]
  wire  _GEN_3548 = fi_sram_idx == 2'h2 ? meta_2_io_valid_r_async & meta_2_io_dirty_r_async : _GEN_3546; // @[Cache.scala 457:38 Cache.scala 459:22]
  wire [5:0] _GEN_3549 = fi_sram_idx == 2'h3 ? fi_line_idx : _GEN_3540; // @[Cache.scala 457:38 Cache.scala 458:28]
  wire  is_dirty = fi_sram_idx == 2'h3 ? meta_3_io_valid_r_async & meta_3_io_dirty_r_async : _GEN_3548; // @[Cache.scala 457:38 Cache.scala 459:22]
  wire  _T_40 = fi_counter_next == 8'h0; // @[Cache.scala 466:33]
  wire [2:0] _GEN_3551 = fi_counter_next == 8'h0 ? 3'h5 : fi_state; // @[Cache.scala 466:42 Cache.scala 467:22 Cache.scala 399:25]
  wire [2:0] _GEN_3554 = _T_12 ? 3'h3 : fi_state; // @[Cache.scala 472:31 Cache.scala 473:20 Cache.scala 399:25]
  wire [2:0] _GEN_3555 = _T_12 ? 3'h4 : fi_state; // @[Cache.scala 477:31 Cache.scala 478:20 Cache.scala 399:25]
  wire [2:0] _GEN_3556 = _T_40 ? 3'h5 : 3'h1; // @[Cache.scala 484:42 Cache.scala 485:22 Cache.scala 487:22]
  wire [7:0] _GEN_3557 = _T_14 ? fi_counter_next : fi_counter; // @[Cache.scala 482:32 Cache.scala 483:22 Cache.scala 402:27]
  wire [2:0] _GEN_3558 = _T_14 ? _GEN_3556 : fi_state; // @[Cache.scala 482:32 Cache.scala 399:25]
  wire [2:0] _GEN_3560 = _T_48 ? 3'h0 : fi_state; // @[Conditional.scala 39:67 Cache.scala 493:18 Cache.scala 399:25]
  wire [7:0] _GEN_3561 = _T_45 ? _GEN_3557 : fi_counter; // @[Conditional.scala 39:67 Cache.scala 402:27]
  wire [2:0] _GEN_3562 = _T_45 ? _GEN_3558 : _GEN_3560; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_3564 = _T_43 ? _GEN_3555 : _GEN_3562; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_3565 = _T_43 ? fi_counter : _GEN_3561; // @[Conditional.scala 39:67 Cache.scala 402:27]
  wire [5:0] _GEN_3570 = _T_35 ? _GEN_3543 : _GEN_3534; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_3571 = _T_35 ? _GEN_3545 : _GEN_3536; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_3572 = _T_35 ? _GEN_3547 : _GEN_3538; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_3573 = _T_35 ? _GEN_3549 : _GEN_3540; // @[Conditional.scala 39:67]
  wire  _io_out_req_valid_T = state == 4'h1; // @[Cache.scala 504:27]
  wire  _io_out_req_valid_T_1 = state == 4'h4; // @[Cache.scala 505:27]
  wire  _io_out_req_valid_T_2 = state == 4'h1 | _io_out_req_valid_T_1; // @[Cache.scala 504:45]
  wire  _io_out_req_valid_T_3 = state == 4'h5; // @[Cache.scala 506:27]
  wire  _io_out_req_valid_T_4 = _io_out_req_valid_T_2 | _io_out_req_valid_T_3; // @[Cache.scala 505:46]
  wire  _io_out_req_valid_T_6 = _io_out_req_valid_T_4 | _fi_update_T; // @[Cache.scala 506:46]
  wire  _io_out_req_valid_T_7 = fi_state == 3'h3; // @[Cache.scala 508:30]
  wire [27:0] io_out_req_bits_addr_hi = s2_addr[31:4]; // @[Cache.scala 512:37]
  wire [31:0] _io_out_req_bits_addr_T = {io_out_req_bits_addr_hi,4'h0}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_3584 = _io_out_req_valid_T ? _io_out_req_bits_addr_T : 32'h0; // @[Cache.scala 511:33 Cache.scala 512:23 Cache.scala 510:21]
  wire [31:0] _io_out_req_bits_addr_T_1 = {1'h1,s2_reg_tag_r,s2_idx,4'h0}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_3585 = _io_out_req_valid_T_1 ? _io_out_req_bits_addr_T_1 : _GEN_3584; // @[Cache.scala 514:34 Cache.scala 517:23]
  wire [31:0] _io_out_req_bits_addr_T_2 = {1'h1,_GEN_3531,fi_line_idx,4'h0}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_3587 = _io_out_req_valid_T_1 ? s2_reg_dat_w[63:0] : 64'h0; // @[Cache.scala 527:34 Cache.scala 528:24 Cache.scala 526:22]
  wire [63:0] _GEN_3588 = _io_out_req_valid_T_3 ? s2_reg_dat_w[127:64] : _GEN_3587; // @[Cache.scala 530:34 Cache.scala 531:24]
  wire [63:0] _GEN_3589 = _fi_update_T ? _GEN_3526[63:0] : _GEN_3588; // @[Cache.scala 533:33 Cache.scala 534:24]
  wire  _io_out_req_bits_wen_T_2 = _io_out_req_valid_T_1 | _io_out_req_valid_T_3; // @[Cache.scala 542:49]
  wire  _io_out_req_bits_wen_T_4 = _io_out_req_bits_wen_T_2 | _fi_update_T; // @[Cache.scala 543:49]
  wire  _io_out_resp_ready_T_1 = state == 4'h6; // @[Cache.scala 549:28]
  wire  _io_out_resp_ready_T_2 = state == 4'h2 | _io_out_resp_ready_T_1; // @[Cache.scala 548:47]
  wire  _io_out_resp_ready_T_3 = fi_state == 3'h4; // @[Cache.scala 550:31]


    assign io_sram4_addr = sram_0_io_addr; 
  assign io_sram4_cen = ~sram_0_io_en; 
  assign io_sram4_wen = ~sram_0_io_wen; 
  assign io_sram4_wdata = sram_0_io_wdata; 
  assign io_sram5_addr = sram_1_io_addr; 
  assign io_sram5_cen = ~sram_1_io_en; 
  assign io_sram5_wen = ~sram_1_io_wen; 
  assign io_sram5_wdata = sram_1_io_wdata; 
  assign io_sram6_addr = sram_2_io_addr; 
  assign io_sram6_cen = ~sram_2_io_en; 
  assign io_sram6_wen = ~sram_2_io_wen; 
  assign io_sram6_wdata = sram_2_io_wdata; 
  assign io_sram7_addr = sram_3_io_addr; 
  assign io_sram7_cen = ~sram_3_io_en; 
  assign io_sram7_wen = ~sram_3_io_wen; 
  assign io_sram7_wdata = sram_3_io_wdata; 

  assign sram_0_io_rdata = io_sram4_rdata;
  assign sram_3_io_rdata = io_sram7_rdata;
  assign sram_2_io_rdata = io_sram6_rdata;
  assign sram_1_io_rdata = io_sram5_rdata;
/*
  ysyx_210340_Sram sram_0 ( // @[Cache.scala 91:22]
    .clock(sram_0_clock),
    .io_en(sram_0_io_en),
    .io_wen(sram_0_io_wen),
    .io_addr(sram_0_io_addr),
    .io_wdata(sram_0_io_wdata),
    .io_rdata(sram_0_io_rdata)
  );
  ysyx_210340_Sram sram_1 ( // @[Cache.scala 91:22]
    .clock(sram_1_clock),
    .io_en(sram_1_io_en),
    .io_wen(sram_1_io_wen),
    .io_addr(sram_1_io_addr),
    .io_wdata(sram_1_io_wdata),
    .io_rdata(sram_1_io_rdata)
  );
  ysyx_210340_Sram sram_2 ( // @[Cache.scala 91:22]
    .clock(sram_2_clock),
    .io_en(sram_2_io_en),
    .io_wen(sram_2_io_wen),
    .io_addr(sram_2_io_addr),
    .io_wdata(sram_2_io_wdata),
    .io_rdata(sram_2_io_rdata)
  );
  ysyx_210340_Sram sram_3 ( // @[Cache.scala 91:22]
    .clock(sram_3_clock),
    .io_en(sram_3_io_en),
    .io_wen(sram_3_io_wen),
    .io_addr(sram_3_io_addr),
    .io_wdata(sram_3_io_wdata),
    .io_rdata(sram_3_io_rdata)
  );
  */
  ysyx_210340_Meta meta_0 ( // @[Cache.scala 99:22]
    .clock(meta_0_clock),
    .reset(meta_0_reset),
    .io_idx(meta_0_io_idx),
    .io_tag_r(meta_0_io_tag_r),
    .io_tag_w(meta_0_io_tag_w),
    .io_tag_wen(meta_0_io_tag_wen),
    .io_dirty_r(meta_0_io_dirty_r),
    .io_dirty_w(meta_0_io_dirty_w),
    .io_dirty_wen(meta_0_io_dirty_wen),
    .io_valid_r(meta_0_io_valid_r),
    .io_invalidate(meta_0_io_invalidate),
    .io_dirty_r_async(meta_0_io_dirty_r_async),
    .io_valid_r_async(meta_0_io_valid_r_async)
  );
  ysyx_210340_Meta meta_1 ( // @[Cache.scala 99:22]
    .clock(meta_1_clock),
    .reset(meta_1_reset),
    .io_idx(meta_1_io_idx),
    .io_tag_r(meta_1_io_tag_r),
    .io_tag_w(meta_1_io_tag_w),
    .io_tag_wen(meta_1_io_tag_wen),
    .io_dirty_r(meta_1_io_dirty_r),
    .io_dirty_w(meta_1_io_dirty_w),
    .io_dirty_wen(meta_1_io_dirty_wen),
    .io_valid_r(meta_1_io_valid_r),
    .io_invalidate(meta_1_io_invalidate),
    .io_dirty_r_async(meta_1_io_dirty_r_async),
    .io_valid_r_async(meta_1_io_valid_r_async)
  );
  ysyx_210340_Meta meta_2 ( // @[Cache.scala 99:22]
    .clock(meta_2_clock),
    .reset(meta_2_reset),
    .io_idx(meta_2_io_idx),
    .io_tag_r(meta_2_io_tag_r),
    .io_tag_w(meta_2_io_tag_w),
    .io_tag_wen(meta_2_io_tag_wen),
    .io_dirty_r(meta_2_io_dirty_r),
    .io_dirty_w(meta_2_io_dirty_w),
    .io_dirty_wen(meta_2_io_dirty_wen),
    .io_valid_r(meta_2_io_valid_r),
    .io_invalidate(meta_2_io_invalidate),
    .io_dirty_r_async(meta_2_io_dirty_r_async),
    .io_valid_r_async(meta_2_io_valid_r_async)
  );
  ysyx_210340_Meta meta_3 ( // @[Cache.scala 99:22]
    .clock(meta_3_clock),
    .reset(meta_3_reset),
    .io_idx(meta_3_io_idx),
    .io_tag_r(meta_3_io_tag_r),
    .io_tag_w(meta_3_io_tag_w),
    .io_tag_wen(meta_3_io_tag_wen),
    .io_dirty_r(meta_3_io_dirty_r),
    .io_dirty_w(meta_3_io_dirty_w),
    .io_dirty_wen(meta_3_io_dirty_wen),
    .io_valid_r(meta_3_io_valid_r),
    .io_invalidate(meta_3_io_invalidate),
    .io_dirty_r_async(meta_3_io_dirty_r_async),
    .io_valid_r_async(meta_3_io_valid_r_async)
  );
  assign io_in_req_ready = fi_ready & ~fi_valid; // @[Cache.scala 275:34]
  assign io_in_resp_valid = s2_hit_real & ~s2_wen & state != 4'h8 | _hit_ready_T; // @[Cache.scala 276:71]
  assign io_in_resp_bits_rdata = _T_2 ? _GEN_228 : _GEN_3295; // @[Conditional.scala 40:58]
  assign io_out_req_valid = _io_out_req_valid_T_6 | _io_out_req_valid_T_7; // @[Cache.scala 507:45]
  assign io_out_req_bits_addr = _fi_update_T ? _io_out_req_bits_addr_T_2 : _GEN_3585; // @[Cache.scala 519:33 Cache.scala 520:23]
  assign io_out_req_bits_aen = _io_out_req_valid_T_2 | _fi_update_T; // @[Cache.scala 523:49]
  assign io_out_req_bits_ren = state == 4'h1; // @[Cache.scala 525:30]
  assign io_out_req_bits_wdata = _io_out_req_valid_T_7 ? _GEN_3526[127:64] : _GEN_3589; // @[Cache.scala 536:33 Cache.scala 537:24]
  assign io_out_req_bits_wlast = _io_out_req_valid_T_3 | _io_out_req_valid_T_7; // @[Cache.scala 540:51]
  assign io_out_req_bits_wen = _io_out_req_bits_wen_T_4 | _io_out_req_valid_T_7; // @[Cache.scala 544:48]
  assign io_out_resp_ready = _io_out_resp_ready_T_2 | _io_out_resp_ready_T_3; // @[Cache.scala 549:47]
  assign dcache_fi_complete_0 = dcache_fi_complete;
  // assign sram_0_clock = clock;
  assign sram_0_io_en = _fi_update_T_1 | _GEN_3489; // @[Cache.scala 437:40 Cache.scala 439:17]
  assign sram_0_io_wen = _T_2 ? _GEN_968 : _GEN_3079; // @[Conditional.scala 40:58]
  assign sram_0_io_addr = _fi_update_T_1 ? fi_line_idx : _GEN_3491; // @[Cache.scala 437:40 Cache.scala 440:19]
  assign sram_0_io_wdata = _T_2 ? _GEN_970 : _GEN_3081; // @[Conditional.scala 40:58]
  // assign sram_1_clock = clock;
  assign sram_1_io_en = _fi_update_T_1 | _GEN_3494; // @[Cache.scala 437:40 Cache.scala 439:17]
  assign sram_1_io_wen = _T_2 ? _GEN_972 : _GEN_3085; // @[Conditional.scala 40:58]
  assign sram_1_io_addr = _fi_update_T_1 ? fi_line_idx : _GEN_3496; // @[Cache.scala 437:40 Cache.scala 440:19]
  assign sram_1_io_wdata = _T_2 ? _GEN_974 : _GEN_3087; // @[Conditional.scala 40:58]
  // assign sram_2_clock = clock;
  assign sram_2_io_en = _fi_update_T_1 | _GEN_3499; // @[Cache.scala 437:40 Cache.scala 439:17]
  assign sram_2_io_wen = _T_2 ? _GEN_976 : _GEN_3091; // @[Conditional.scala 40:58]
  assign sram_2_io_addr = _fi_update_T_1 ? fi_line_idx : _GEN_3501; // @[Cache.scala 437:40 Cache.scala 440:19]
  assign sram_2_io_wdata = _T_2 ? _GEN_978 : _GEN_3093; // @[Conditional.scala 40:58]
  // assign sram_3_clock = clock;
  assign sram_3_io_en = _fi_update_T_1 | _GEN_3504; // @[Cache.scala 437:40 Cache.scala 439:17]
  assign sram_3_io_wen = _T_2 ? _GEN_980 : _GEN_3097; // @[Conditional.scala 40:58]
  assign sram_3_io_addr = _fi_update_T_1 ? fi_line_idx : _GEN_3506; // @[Cache.scala 437:40 Cache.scala 440:19]
  assign sram_3_io_wdata = _T_2 ? _GEN_982 : _GEN_3099; // @[Conditional.scala 40:58]
  assign meta_0_clock = clock;
  assign meta_0_reset = reset;
  assign meta_0_io_idx = _T_34 ? _GEN_3534 : _GEN_3570; // @[Conditional.scala 40:58]
  assign meta_0_io_tag_w = _T_2 ? 21'h0 : _GEN_3082; // @[Conditional.scala 40:58 Cache.scala 116:16]
  assign meta_0_io_tag_wen = _T_2 ? 1'h0 : _GEN_3079; // @[Conditional.scala 40:58 Cache.scala 117:18]
  assign meta_0_io_dirty_w = _T_2 ? _GEN_968 : _GEN_3083; // @[Conditional.scala 40:58]
  assign meta_0_io_dirty_wen = _T_2 ? _GEN_968 : _GEN_3079; // @[Conditional.scala 40:58]
  assign meta_0_io_invalidate = _T_34 ? 1'h0 : _GEN_3576; // @[Conditional.scala 40:58]
  assign meta_1_clock = clock;
  assign meta_1_reset = reset;
  assign meta_1_io_idx = _T_34 ? _GEN_3536 : _GEN_3571; // @[Conditional.scala 40:58]
  assign meta_1_io_tag_w = _T_2 ? 21'h0 : _GEN_3088; // @[Conditional.scala 40:58 Cache.scala 116:16]
  assign meta_1_io_tag_wen = _T_2 ? 1'h0 : _GEN_3085; // @[Conditional.scala 40:58 Cache.scala 117:18]
  assign meta_1_io_dirty_w = _T_2 ? _GEN_972 : _GEN_3089; // @[Conditional.scala 40:58]
  assign meta_1_io_dirty_wen = _T_2 ? _GEN_972 : _GEN_3085; // @[Conditional.scala 40:58]
  assign meta_1_io_invalidate = _T_34 ? 1'h0 : _GEN_3576; // @[Conditional.scala 40:58]
  assign meta_2_clock = clock;
  assign meta_2_reset = reset;
  assign meta_2_io_idx = _T_34 ? _GEN_3538 : _GEN_3572; // @[Conditional.scala 40:58]
  assign meta_2_io_tag_w = _T_2 ? 21'h0 : _GEN_3094; // @[Conditional.scala 40:58 Cache.scala 116:16]
  assign meta_2_io_tag_wen = _T_2 ? 1'h0 : _GEN_3091; // @[Conditional.scala 40:58 Cache.scala 117:18]
  assign meta_2_io_dirty_w = _T_2 ? _GEN_976 : _GEN_3095; // @[Conditional.scala 40:58]
  assign meta_2_io_dirty_wen = _T_2 ? _GEN_976 : _GEN_3091; // @[Conditional.scala 40:58]
  assign meta_2_io_invalidate = _T_34 ? 1'h0 : _GEN_3576; // @[Conditional.scala 40:58]
  assign meta_3_clock = clock;
  assign meta_3_reset = reset;
  assign meta_3_io_idx = _T_34 ? _GEN_3540 : _GEN_3573; // @[Conditional.scala 40:58]
  assign meta_3_io_tag_w = _T_2 ? 21'h0 : _GEN_3100; // @[Conditional.scala 40:58 Cache.scala 116:16]
  assign meta_3_io_tag_wen = _T_2 ? 1'h0 : _GEN_3097; // @[Conditional.scala 40:58 Cache.scala 117:18]
  assign meta_3_io_dirty_w = _T_2 ? _GEN_980 : _GEN_3101; // @[Conditional.scala 40:58]
  assign meta_3_io_dirty_wen = _T_2 ? _GEN_980 : _GEN_3097; // @[Conditional.scala 40:58]
  assign meta_3_io_invalidate = _T_34 ? 1'h0 : _GEN_3576; // @[Conditional.scala 40:58]
  always @(posedge clock) begin
    if (reset) begin // @[Cache.scala 131:22]
      plru0_0 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_0 <= _GEN_229;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_0 <= _GEN_2660;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_1 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_1 <= _GEN_230;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_1 <= _GEN_2661;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_2 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_2 <= _GEN_231;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_2 <= _GEN_2662;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_3 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_3 <= _GEN_232;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_3 <= _GEN_2663;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_4 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_4 <= _GEN_233;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_4 <= _GEN_2664;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_5 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_5 <= _GEN_234;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_5 <= _GEN_2665;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_6 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_6 <= _GEN_235;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_6 <= _GEN_2666;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_7 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_7 <= _GEN_236;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_7 <= _GEN_2667;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_8 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_8 <= _GEN_237;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_8 <= _GEN_2668;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_9 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_9 <= _GEN_238;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_9 <= _GEN_2669;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_10 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_10 <= _GEN_239;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_10 <= _GEN_2670;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_11 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_11 <= _GEN_240;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_11 <= _GEN_2671;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_12 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_12 <= _GEN_241;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_12 <= _GEN_2672;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_13 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_13 <= _GEN_242;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_13 <= _GEN_2673;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_14 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_14 <= _GEN_243;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_14 <= _GEN_2674;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_15 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_15 <= _GEN_244;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_15 <= _GEN_2675;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_16 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_16 <= _GEN_245;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_16 <= _GEN_2676;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_17 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_17 <= _GEN_246;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_17 <= _GEN_2677;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_18 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_18 <= _GEN_247;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_18 <= _GEN_2678;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_19 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_19 <= _GEN_248;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_19 <= _GEN_2679;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_20 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_20 <= _GEN_249;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_20 <= _GEN_2680;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_21 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_21 <= _GEN_250;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_21 <= _GEN_2681;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_22 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_22 <= _GEN_251;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_22 <= _GEN_2682;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_23 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_23 <= _GEN_252;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_23 <= _GEN_2683;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_24 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_24 <= _GEN_253;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_24 <= _GEN_2684;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_25 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_25 <= _GEN_254;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_25 <= _GEN_2685;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_26 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_26 <= _GEN_255;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_26 <= _GEN_2686;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_27 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_27 <= _GEN_256;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_27 <= _GEN_2687;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_28 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_28 <= _GEN_257;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_28 <= _GEN_2688;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_29 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_29 <= _GEN_258;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_29 <= _GEN_2689;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_30 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_30 <= _GEN_259;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_30 <= _GEN_2690;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_31 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_31 <= _GEN_260;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_31 <= _GEN_2691;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_32 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_32 <= _GEN_261;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_32 <= _GEN_2692;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_33 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_33 <= _GEN_262;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_33 <= _GEN_2693;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_34 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_34 <= _GEN_263;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_34 <= _GEN_2694;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_35 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_35 <= _GEN_264;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_35 <= _GEN_2695;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_36 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_36 <= _GEN_265;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_36 <= _GEN_2696;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_37 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_37 <= _GEN_266;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_37 <= _GEN_2697;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_38 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_38 <= _GEN_267;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_38 <= _GEN_2698;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_39 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_39 <= _GEN_268;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_39 <= _GEN_2699;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_40 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_40 <= _GEN_269;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_40 <= _GEN_2700;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_41 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_41 <= _GEN_270;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_41 <= _GEN_2701;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_42 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_42 <= _GEN_271;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_42 <= _GEN_2702;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_43 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_43 <= _GEN_272;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_43 <= _GEN_2703;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_44 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_44 <= _GEN_273;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_44 <= _GEN_2704;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_45 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_45 <= _GEN_274;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_45 <= _GEN_2705;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_46 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_46 <= _GEN_275;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_46 <= _GEN_2706;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_47 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_47 <= _GEN_276;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_47 <= _GEN_2707;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_48 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_48 <= _GEN_277;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_48 <= _GEN_2708;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_49 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_49 <= _GEN_278;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_49 <= _GEN_2709;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_50 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_50 <= _GEN_279;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_50 <= _GEN_2710;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_51 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_51 <= _GEN_280;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_51 <= _GEN_2711;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_52 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_52 <= _GEN_281;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_52 <= _GEN_2712;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_53 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_53 <= _GEN_282;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_53 <= _GEN_2713;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_54 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_54 <= _GEN_283;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_54 <= _GEN_2714;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_55 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_55 <= _GEN_284;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_55 <= _GEN_2715;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_56 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_56 <= _GEN_285;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_56 <= _GEN_2716;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_57 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_57 <= _GEN_286;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_57 <= _GEN_2717;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_58 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_58 <= _GEN_287;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_58 <= _GEN_2718;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_59 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_59 <= _GEN_288;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_59 <= _GEN_2719;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_60 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_60 <= _GEN_289;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_60 <= _GEN_2720;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_61 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_61 <= _GEN_290;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_61 <= _GEN_2721;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_62 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_62 <= _GEN_291;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_62 <= _GEN_2722;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru0_63 <= 1'h0; // @[Cache.scala 131:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru0_63 <= _GEN_292;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru0_63 <= _GEN_2723;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_0 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_0 <= _GEN_421;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_0 <= _GEN_2724;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_1 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_1 <= _GEN_422;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_1 <= _GEN_2725;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_2 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_2 <= _GEN_423;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_2 <= _GEN_2726;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_3 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_3 <= _GEN_424;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_3 <= _GEN_2727;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_4 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_4 <= _GEN_425;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_4 <= _GEN_2728;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_5 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_5 <= _GEN_426;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_5 <= _GEN_2729;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_6 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_6 <= _GEN_427;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_6 <= _GEN_2730;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_7 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_7 <= _GEN_428;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_7 <= _GEN_2731;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_8 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_8 <= _GEN_429;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_8 <= _GEN_2732;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_9 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_9 <= _GEN_430;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_9 <= _GEN_2733;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_10 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_10 <= _GEN_431;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_10 <= _GEN_2734;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_11 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_11 <= _GEN_432;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_11 <= _GEN_2735;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_12 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_12 <= _GEN_433;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_12 <= _GEN_2736;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_13 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_13 <= _GEN_434;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_13 <= _GEN_2737;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_14 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_14 <= _GEN_435;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_14 <= _GEN_2738;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_15 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_15 <= _GEN_436;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_15 <= _GEN_2739;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_16 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_16 <= _GEN_437;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_16 <= _GEN_2740;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_17 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_17 <= _GEN_438;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_17 <= _GEN_2741;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_18 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_18 <= _GEN_439;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_18 <= _GEN_2742;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_19 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_19 <= _GEN_440;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_19 <= _GEN_2743;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_20 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_20 <= _GEN_441;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_20 <= _GEN_2744;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_21 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_21 <= _GEN_442;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_21 <= _GEN_2745;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_22 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_22 <= _GEN_443;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_22 <= _GEN_2746;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_23 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_23 <= _GEN_444;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_23 <= _GEN_2747;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_24 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_24 <= _GEN_445;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_24 <= _GEN_2748;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_25 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_25 <= _GEN_446;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_25 <= _GEN_2749;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_26 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_26 <= _GEN_447;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_26 <= _GEN_2750;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_27 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_27 <= _GEN_448;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_27 <= _GEN_2751;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_28 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_28 <= _GEN_449;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_28 <= _GEN_2752;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_29 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_29 <= _GEN_450;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_29 <= _GEN_2753;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_30 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_30 <= _GEN_451;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_30 <= _GEN_2754;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_31 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_31 <= _GEN_452;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_31 <= _GEN_2755;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_32 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_32 <= _GEN_453;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_32 <= _GEN_2756;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_33 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_33 <= _GEN_454;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_33 <= _GEN_2757;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_34 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_34 <= _GEN_455;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_34 <= _GEN_2758;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_35 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_35 <= _GEN_456;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_35 <= _GEN_2759;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_36 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_36 <= _GEN_457;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_36 <= _GEN_2760;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_37 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_37 <= _GEN_458;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_37 <= _GEN_2761;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_38 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_38 <= _GEN_459;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_38 <= _GEN_2762;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_39 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_39 <= _GEN_460;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_39 <= _GEN_2763;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_40 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_40 <= _GEN_461;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_40 <= _GEN_2764;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_41 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_41 <= _GEN_462;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_41 <= _GEN_2765;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_42 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_42 <= _GEN_463;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_42 <= _GEN_2766;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_43 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_43 <= _GEN_464;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_43 <= _GEN_2767;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_44 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_44 <= _GEN_465;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_44 <= _GEN_2768;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_45 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_45 <= _GEN_466;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_45 <= _GEN_2769;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_46 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_46 <= _GEN_467;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_46 <= _GEN_2770;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_47 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_47 <= _GEN_468;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_47 <= _GEN_2771;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_48 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_48 <= _GEN_469;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_48 <= _GEN_2772;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_49 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_49 <= _GEN_470;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_49 <= _GEN_2773;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_50 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_50 <= _GEN_471;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_50 <= _GEN_2774;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_51 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_51 <= _GEN_472;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_51 <= _GEN_2775;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_52 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_52 <= _GEN_473;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_52 <= _GEN_2776;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_53 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_53 <= _GEN_474;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_53 <= _GEN_2777;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_54 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_54 <= _GEN_475;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_54 <= _GEN_2778;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_55 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_55 <= _GEN_476;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_55 <= _GEN_2779;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_56 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_56 <= _GEN_477;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_56 <= _GEN_2780;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_57 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_57 <= _GEN_478;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_57 <= _GEN_2781;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_58 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_58 <= _GEN_479;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_58 <= _GEN_2782;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_59 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_59 <= _GEN_480;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_59 <= _GEN_2783;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_60 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_60 <= _GEN_481;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_60 <= _GEN_2784;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_61 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_61 <= _GEN_482;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_61 <= _GEN_2785;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_62 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_62 <= _GEN_483;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_62 <= _GEN_2786;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru1_63 <= 1'h0; // @[Cache.scala 133:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru1_63 <= _GEN_484;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru1_63 <= _GEN_2787;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_0 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_0 <= _GEN_485;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_0 <= _GEN_2788;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_1 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_1 <= _GEN_486;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_1 <= _GEN_2789;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_2 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_2 <= _GEN_487;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_2 <= _GEN_2790;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_3 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_3 <= _GEN_488;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_3 <= _GEN_2791;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_4 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_4 <= _GEN_489;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_4 <= _GEN_2792;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_5 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_5 <= _GEN_490;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_5 <= _GEN_2793;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_6 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_6 <= _GEN_491;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_6 <= _GEN_2794;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_7 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_7 <= _GEN_492;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_7 <= _GEN_2795;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_8 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_8 <= _GEN_493;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_8 <= _GEN_2796;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_9 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_9 <= _GEN_494;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_9 <= _GEN_2797;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_10 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_10 <= _GEN_495;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_10 <= _GEN_2798;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_11 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_11 <= _GEN_496;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_11 <= _GEN_2799;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_12 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_12 <= _GEN_497;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_12 <= _GEN_2800;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_13 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_13 <= _GEN_498;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_13 <= _GEN_2801;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_14 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_14 <= _GEN_499;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_14 <= _GEN_2802;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_15 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_15 <= _GEN_500;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_15 <= _GEN_2803;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_16 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_16 <= _GEN_501;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_16 <= _GEN_2804;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_17 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_17 <= _GEN_502;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_17 <= _GEN_2805;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_18 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_18 <= _GEN_503;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_18 <= _GEN_2806;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_19 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_19 <= _GEN_504;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_19 <= _GEN_2807;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_20 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_20 <= _GEN_505;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_20 <= _GEN_2808;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_21 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_21 <= _GEN_506;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_21 <= _GEN_2809;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_22 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_22 <= _GEN_507;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_22 <= _GEN_2810;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_23 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_23 <= _GEN_508;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_23 <= _GEN_2811;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_24 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_24 <= _GEN_509;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_24 <= _GEN_2812;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_25 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_25 <= _GEN_510;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_25 <= _GEN_2813;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_26 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_26 <= _GEN_511;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_26 <= _GEN_2814;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_27 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_27 <= _GEN_512;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_27 <= _GEN_2815;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_28 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_28 <= _GEN_513;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_28 <= _GEN_2816;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_29 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_29 <= _GEN_514;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_29 <= _GEN_2817;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_30 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_30 <= _GEN_515;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_30 <= _GEN_2818;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_31 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_31 <= _GEN_516;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_31 <= _GEN_2819;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_32 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_32 <= _GEN_517;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_32 <= _GEN_2820;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_33 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_33 <= _GEN_518;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_33 <= _GEN_2821;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_34 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_34 <= _GEN_519;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_34 <= _GEN_2822;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_35 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_35 <= _GEN_520;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_35 <= _GEN_2823;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_36 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_36 <= _GEN_521;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_36 <= _GEN_2824;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_37 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_37 <= _GEN_522;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_37 <= _GEN_2825;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_38 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_38 <= _GEN_523;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_38 <= _GEN_2826;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_39 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_39 <= _GEN_524;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_39 <= _GEN_2827;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_40 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_40 <= _GEN_525;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_40 <= _GEN_2828;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_41 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_41 <= _GEN_526;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_41 <= _GEN_2829;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_42 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_42 <= _GEN_527;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_42 <= _GEN_2830;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_43 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_43 <= _GEN_528;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_43 <= _GEN_2831;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_44 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_44 <= _GEN_529;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_44 <= _GEN_2832;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_45 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_45 <= _GEN_530;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_45 <= _GEN_2833;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_46 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_46 <= _GEN_531;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_46 <= _GEN_2834;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_47 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_47 <= _GEN_532;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_47 <= _GEN_2835;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_48 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_48 <= _GEN_533;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_48 <= _GEN_2836;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_49 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_49 <= _GEN_534;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_49 <= _GEN_2837;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_50 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_50 <= _GEN_535;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_50 <= _GEN_2838;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_51 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_51 <= _GEN_536;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_51 <= _GEN_2839;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_52 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_52 <= _GEN_537;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_52 <= _GEN_2840;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_53 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_53 <= _GEN_538;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_53 <= _GEN_2841;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_54 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_54 <= _GEN_539;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_54 <= _GEN_2842;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_55 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_55 <= _GEN_540;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_55 <= _GEN_2843;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_56 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_56 <= _GEN_541;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_56 <= _GEN_2844;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_57 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_57 <= _GEN_542;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_57 <= _GEN_2845;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_58 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_58 <= _GEN_543;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_58 <= _GEN_2846;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_59 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_59 <= _GEN_544;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_59 <= _GEN_2847;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_60 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_60 <= _GEN_545;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_60 <= _GEN_2848;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_61 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_61 <= _GEN_546;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_61 <= _GEN_2849;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_62 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_62 <= _GEN_547;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_62 <= _GEN_2850;
      end
    end
    if (reset) begin // @[Cache.scala 135:22]
      plru2_63 <= 1'h0; // @[Cache.scala 135:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (REG_2) begin // @[Cache.scala 289:37]
        if (s2_hit) begin // @[Cache.scala 290:23]
          plru2_63 <= _GEN_548;
        end
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_13)) begin // @[Conditional.scala 39:67]
        plru2_63 <= _GEN_2851;
      end
    end
    s2_hit_real_REG <= (hit_ready | _hit_ready_T) & io_in_resp_ready | invalid_ready; // @[Cache.scala 270:66]
    if (reset) begin // @[Cache.scala 209:25]
      s2_addr <= 32'h0; // @[Cache.scala 209:25]
    end else if (fi_ready) begin // @[Cache.scala 238:24]
      s2_addr <= io_in_req_bits_addr; // @[Cache.scala 240:14]
    end
    if (reset) begin // @[Cache.scala 231:27]
      s2_reg_hit <= 1'h0; // @[Cache.scala 231:27]
    end else if (!(fi_ready)) begin // @[Cache.scala 238:24]
      if (~fi_ready & REG) begin // @[Cache.scala 244:58]
        s2_reg_hit <= s2_hit; // @[Cache.scala 247:18]
      end
    end
    if (reset) begin // @[Cache.scala 213:25]
      s2_wen <= 1'h0; // @[Cache.scala 213:25]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      s2_wen <= _GEN_27;
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      s2_wen <= _GEN_27;
    end else if (_T_13) begin // @[Conditional.scala 39:67]
      s2_wen <= _GEN_27;
    end else begin
      s2_wen <= _GEN_2852;
    end
    if (reset) begin // @[Cache.scala 207:22]
      state <= 4'h8; // @[Cache.scala 207:22]
    end else if (fi_fire) begin // @[Cache.scala 411:18]
      state <= 4'h8; // @[Cache.scala 412:11]
    end else if (fi_ready) begin // @[Cache.scala 381:24]
      if (io_in_req_valid) begin // @[Cache.scala 382:17]
        state <= 4'h0;
      end else begin
        state <= 4'h8;
      end
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      state <= _GEN_983;
    end else begin
      state <= _GEN_3075;
    end
    if (reset) begin // @[ID.scala 18:20]
      fi_valid <= 1'h0; // @[ID.scala 18:20]
    end else if (dcache_fi_complete) begin // @[ID.scala 25:19]
      fi_valid <= 1'h0; // @[ID.scala 25:23]
    end else begin
      fi_valid <= _GEN_0;
    end
    if (reset) begin // @[Cache.scala 399:25]
      fi_state <= 3'h0; // @[Cache.scala 399:25]
    end else if (_T_34) begin // @[Conditional.scala 40:58]
      if (fi_fire) begin // @[Cache.scala 449:24]
        fi_state <= 3'h1; // @[Cache.scala 451:20]
      end
    end else if (_T_35) begin // @[Conditional.scala 39:67]
      if (is_dirty) begin // @[Cache.scala 462:25]
        fi_state <= 3'h2; // @[Cache.scala 463:20]
      end else begin
        fi_state <= _GEN_3551;
      end
    end else if (_T_41) begin // @[Conditional.scala 39:67]
      fi_state <= _GEN_3554;
    end else begin
      fi_state <= _GEN_3564;
    end
    if (reset) begin // @[Cache.scala 214:25]
      s2_wdata <= 64'h0; // @[Cache.scala 214:25]
    end else if (fi_ready) begin // @[Cache.scala 238:24]
      s2_wdata <= io_in_req_bits_wdata; // @[Cache.scala 242:14]
    end
    if (reset) begin // @[Cache.scala 215:25]
      s2_wmask <= 8'h0; // @[Cache.scala 215:25]
    end else if (fi_ready) begin // @[Cache.scala 238:24]
      s2_wmask <= io_in_req_bits_wmask; // @[Cache.scala 243:14]
    end
    if (reset) begin // @[Cache.scala 233:29]
      s2_reg_rdata <= 128'h0; // @[Cache.scala 233:29]
    end else if (!(fi_ready)) begin // @[Cache.scala 238:24]
      if (~fi_ready & REG) begin // @[Cache.scala 244:58]
        if (2'h3 == s2_way) begin // @[Cache.scala 249:18]
          s2_reg_rdata <= sram_out_3; // @[Cache.scala 249:18]
        end else begin
          s2_reg_rdata <= _GEN_6;
        end
      end
    end
    if (reset) begin // @[Cache.scala 234:29]
      s2_reg_dirty <= 1'h0; // @[Cache.scala 234:29]
    end else if (!(fi_ready)) begin // @[Cache.scala 238:24]
      if (~fi_ready & REG) begin // @[Cache.scala 244:58]
        if (2'h3 == replace_way) begin // @[Cache.scala 250:18]
          s2_reg_dirty <= dirty_out_3; // @[Cache.scala 250:18]
        end else begin
          s2_reg_dirty <= _GEN_10;
        end
      end
    end
    if (reset) begin // @[Cache.scala 235:29]
      s2_reg_tag_r <= 21'h0; // @[Cache.scala 235:29]
    end else if (!(fi_ready)) begin // @[Cache.scala 238:24]
      if (~fi_ready & REG) begin // @[Cache.scala 244:58]
        if (2'h3 == replace_way) begin // @[Cache.scala 251:18]
          s2_reg_tag_r <= tag_out_3; // @[Cache.scala 251:18]
        end else begin
          s2_reg_tag_r <= _GEN_14;
        end
      end
    end
    if (reset) begin // @[Cache.scala 236:29]
      s2_reg_dat_w <= 128'h0; // @[Cache.scala 236:29]
    end else if (!(fi_ready)) begin // @[Cache.scala 238:24]
      if (~fi_ready & REG) begin // @[Cache.scala 244:58]
        if (2'h3 == replace_way) begin // @[Cache.scala 252:18]
          s2_reg_dat_w <= sram_out_3; // @[Cache.scala 252:18]
        end else begin
          s2_reg_dat_w <= _GEN_18;
        end
      end
    end
    REG <= (hit_ready | _hit_ready_T) & io_in_resp_ready | invalid_ready; // @[Cache.scala 270:66]
    if (reset) begin // @[Cache.scala 258:23]
      wdata1 <= 64'h0; // @[Cache.scala 258:23]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (!(_T_11)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          wdata1 <= _GEN_988;
        end
      end
    end
    if (reset) begin // @[Cache.scala 259:23]
      wdata2 <= 64'h0; // @[Cache.scala 259:23]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (!(_T_11)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          wdata2 <= _GEN_989;
        end
      end
    end
    REG_1 <= (hit_ready | _hit_ready_T) & io_in_resp_ready | invalid_ready; // @[Cache.scala 270:66]
    REG_2 <= (hit_ready | _hit_ready_T) & io_in_resp_ready | invalid_ready; // @[Cache.scala 270:66]
    if (s2_offs) begin // @[Cache.scala 374:40]
      io_in_resp_bits_rdata_REG <= wdata2;
    end else begin
      io_in_resp_bits_rdata_REG <= wdata1;
    end
    if (reset) begin // @[Cache.scala 402:27]
      fi_counter <= 8'h0; // @[Cache.scala 402:27]
    end else if (_T_34) begin // @[Conditional.scala 40:58]
      if (fi_fire) begin // @[Cache.scala 449:24]
        fi_counter <= 8'h0; // @[Cache.scala 450:22]
      end
    end else if (_T_35) begin // @[Conditional.scala 39:67]
      if (!(is_dirty)) begin // @[Cache.scala 462:25]
        fi_counter <= fi_counter_next; // @[Cache.scala 465:22]
      end
    end else if (!(_T_41)) begin // @[Conditional.scala 39:67]
      fi_counter <= _GEN_3565;
    end
    fi_update_REG <= fi_state == 3'h1; // @[Cache.scala 407:65]
    if (reset) begin // @[Reg.scala 27:20]
      fi_wdata_r <= 128'h0; // @[Reg.scala 27:20]
    end else if (fi_update) begin // @[Reg.scala 28:19]
      if (2'h3 == fi_sram_idx) begin // @[Reg.scala 28:23]
        fi_wdata_r <= sram_out_3; // @[Reg.scala 28:23]
      end else if (2'h2 == fi_sram_idx) begin // @[Reg.scala 28:23]
        fi_wdata_r <= sram_out_2; // @[Reg.scala 28:23]
      end else begin
        fi_wdata_r <= _GEN_3523;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      fi_tag_r <= 21'h0; // @[Reg.scala 27:20]
    end else if (fi_update) begin // @[Reg.scala 28:19]
      if (2'h3 == fi_sram_idx) begin // @[Reg.scala 28:23]
        fi_tag_r <= tag_out_3; // @[Reg.scala 28:23]
      end else if (2'h2 == fi_sram_idx) begin // @[Reg.scala 28:23]
        fi_tag_r <= tag_out_2; // @[Reg.scala 28:23]
      end else begin
        fi_tag_r <= _GEN_3528;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  plru0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  plru0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  plru0_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  plru0_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  plru0_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  plru0_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  plru0_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  plru0_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  plru0_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  plru0_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  plru0_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  plru0_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  plru0_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  plru0_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  plru0_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  plru0_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  plru0_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  plru0_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  plru0_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  plru0_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  plru0_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  plru0_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  plru0_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  plru0_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  plru0_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  plru0_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  plru0_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  plru0_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  plru0_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  plru0_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  plru0_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  plru0_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  plru0_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  plru0_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  plru0_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  plru0_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  plru0_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  plru0_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  plru0_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  plru0_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  plru0_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  plru0_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  plru0_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  plru0_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  plru0_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  plru0_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  plru0_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  plru0_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  plru0_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  plru0_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  plru0_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  plru0_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  plru0_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  plru0_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  plru0_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  plru0_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  plru0_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  plru0_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  plru0_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  plru0_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  plru0_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  plru0_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  plru0_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  plru0_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  plru1_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  plru1_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  plru1_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  plru1_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  plru1_4 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  plru1_5 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  plru1_6 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  plru1_7 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  plru1_8 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  plru1_9 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  plru1_10 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  plru1_11 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  plru1_12 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  plru1_13 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  plru1_14 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  plru1_15 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  plru1_16 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  plru1_17 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  plru1_18 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  plru1_19 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  plru1_20 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  plru1_21 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  plru1_22 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  plru1_23 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  plru1_24 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  plru1_25 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  plru1_26 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  plru1_27 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  plru1_28 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  plru1_29 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  plru1_30 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  plru1_31 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  plru1_32 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  plru1_33 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  plru1_34 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  plru1_35 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  plru1_36 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  plru1_37 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  plru1_38 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  plru1_39 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  plru1_40 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  plru1_41 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  plru1_42 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  plru1_43 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  plru1_44 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  plru1_45 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  plru1_46 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  plru1_47 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  plru1_48 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  plru1_49 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  plru1_50 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  plru1_51 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  plru1_52 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  plru1_53 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  plru1_54 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  plru1_55 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  plru1_56 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  plru1_57 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  plru1_58 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  plru1_59 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  plru1_60 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  plru1_61 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  plru1_62 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  plru1_63 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  plru2_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  plru2_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  plru2_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  plru2_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  plru2_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  plru2_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  plru2_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  plru2_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  plru2_8 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  plru2_9 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  plru2_10 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  plru2_11 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  plru2_12 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  plru2_13 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  plru2_14 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  plru2_15 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  plru2_16 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  plru2_17 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  plru2_18 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  plru2_19 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  plru2_20 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  plru2_21 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  plru2_22 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  plru2_23 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  plru2_24 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  plru2_25 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  plru2_26 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  plru2_27 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  plru2_28 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  plru2_29 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  plru2_30 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  plru2_31 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  plru2_32 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  plru2_33 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  plru2_34 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  plru2_35 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  plru2_36 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  plru2_37 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  plru2_38 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  plru2_39 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  plru2_40 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  plru2_41 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  plru2_42 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  plru2_43 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  plru2_44 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  plru2_45 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  plru2_46 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  plru2_47 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  plru2_48 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  plru2_49 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  plru2_50 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  plru2_51 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  plru2_52 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  plru2_53 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  plru2_54 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  plru2_55 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  plru2_56 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  plru2_57 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  plru2_58 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  plru2_59 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  plru2_60 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  plru2_61 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  plru2_62 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  plru2_63 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  s2_hit_real_REG = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  s2_addr = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  s2_reg_hit = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  s2_wen = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  state = _RAND_196[3:0];
  _RAND_197 = {1{`RANDOM}};
  fi_valid = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  fi_state = _RAND_198[2:0];
  _RAND_199 = {2{`RANDOM}};
  s2_wdata = _RAND_199[63:0];
  _RAND_200 = {1{`RANDOM}};
  s2_wmask = _RAND_200[7:0];
  _RAND_201 = {4{`RANDOM}};
  s2_reg_rdata = _RAND_201[127:0];
  _RAND_202 = {1{`RANDOM}};
  s2_reg_dirty = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  s2_reg_tag_r = _RAND_203[20:0];
  _RAND_204 = {4{`RANDOM}};
  s2_reg_dat_w = _RAND_204[127:0];
  _RAND_205 = {1{`RANDOM}};
  REG = _RAND_205[0:0];
  _RAND_206 = {2{`RANDOM}};
  wdata1 = _RAND_206[63:0];
  _RAND_207 = {2{`RANDOM}};
  wdata2 = _RAND_207[63:0];
  _RAND_208 = {1{`RANDOM}};
  REG_1 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  REG_2 = _RAND_209[0:0];
  _RAND_210 = {2{`RANDOM}};
  io_in_resp_bits_rdata_REG = _RAND_210[63:0];
  _RAND_211 = {1{`RANDOM}};
  fi_counter = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  fi_update_REG = _RAND_212[0:0];
  _RAND_213 = {4{`RANDOM}};
  fi_wdata_r = _RAND_213[127:0];
  _RAND_214 = {1{`RANDOM}};
  fi_tag_r = _RAND_214[20:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210340_Uncache_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input         io_in_req_bits_ren,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input  [1:0]  io_in_req_bits_size,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output        io_out_req_bits_ren,
  output [63:0] io_out_req_bits_wdata,
  output [7:0]  io_out_req_bits_wmask,
  output        io_out_req_bits_wen,
  output [1:0]  io_out_req_bits_size,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[Uncache.scala 18:22]
  reg [31:0] addr; // @[Uncache.scala 21:22]
  reg  ren; // @[Uncache.scala 22:22]
  reg [63:0] wdata; // @[Uncache.scala 23:22]
  reg [7:0] wmask; // @[Uncache.scala 24:22]
  reg  wen; // @[Uncache.scala 25:22]
  reg [1:0] size; // @[Uncache.scala 26:22]
  reg [63:0] rdata_1; // @[Uncache.scala 29:24]
  reg [63:0] rdata_2; // @[Uncache.scala 30:24]
  wire  req_split = size == 2'h3; // @[Uncache.scala 34:22]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_2 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_5 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _state_T = req_split ? 3'h3 : 3'h5; // @[Uncache.scala 59:21]
  wire [63:0] _GEN_10 = _T_5 ? io_out_resp_bits_rdata : rdata_1; // @[Uncache.scala 57:30 Uncache.scala 58:17 Uncache.scala 29:24]
  wire [2:0] _GEN_11 = _T_5 ? _state_T : state; // @[Uncache.scala 57:30 Uncache.scala 59:15 Uncache.scala 18:22]
  wire  _T_6 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_12 = _T_3 ? 3'h4 : state; // @[Uncache.scala 63:29 Uncache.scala 64:15 Uncache.scala 18:22]
  wire  _T_8 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire [63:0] _GEN_13 = _T_5 ? io_out_resp_bits_rdata : rdata_2; // @[Uncache.scala 68:30 Uncache.scala 69:17 Uncache.scala 30:24]
  wire [2:0] _GEN_14 = _T_5 ? 3'h5 : state; // @[Uncache.scala 68:30 Uncache.scala 70:15 Uncache.scala 18:22]
  wire  _T_10 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_11 = io_in_resp_ready & io_in_resp_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_15 = _T_11 ? 3'h0 : state; // @[Uncache.scala 74:29 Uncache.scala 75:15 Uncache.scala 18:22]
  wire [2:0] _GEN_16 = _T_10 ? _GEN_15 : state; // @[Conditional.scala 39:67 Uncache.scala 18:22]
  wire [63:0] _GEN_17 = _T_8 ? _GEN_13 : rdata_2; // @[Conditional.scala 39:67 Uncache.scala 30:24]
  wire [2:0] _GEN_18 = _T_8 ? _GEN_14 : _GEN_16; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_19 = _T_6 ? _GEN_12 : _GEN_18; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_20 = _T_6 ? rdata_2 : _GEN_17; // @[Conditional.scala 39:67 Uncache.scala 30:24]
  wire  _io_out_req_valid_T_1 = state == 3'h3; // @[Uncache.scala 81:55]
  wire [31:0] io_in_resp_bits_rdata_hi = rdata_2[31:0]; // @[Uncache.scala 91:53]
  wire [31:0] io_in_resp_bits_rdata_lo = rdata_1[31:0]; // @[Uncache.scala 91:68]
  wire [63:0] _io_in_resp_bits_rdata_T = {io_in_resp_bits_rdata_hi,io_in_resp_bits_rdata_lo}; // @[Cat.scala 30:58]
  wire [31:0] _io_out_req_bits_addr_T_3 = addr + 32'h4; // @[Uncache.scala 94:70]
  assign io_in_req_ready = state == 3'h0; // @[Uncache.scala 80:34]
  assign io_in_resp_valid = state == 3'h5; // @[Uncache.scala 90:34]
  assign io_in_resp_bits_rdata = req_split ? _io_in_resp_bits_rdata_T : rdata_1; // @[Uncache.scala 91:30]
  assign io_out_req_valid = state == 3'h1 | state == 3'h3; // @[Uncache.scala 81:46]
  assign io_out_req_bits_addr = req_split & _io_out_req_valid_T_1 ? _io_out_req_bits_addr_T_3 : addr; // @[Uncache.scala 94:30]
  assign io_out_req_bits_ren = ren; // @[Uncache.scala 84:24]
  assign io_out_req_bits_wdata = wdata; // @[Uncache.scala 95:24]
  assign io_out_req_bits_wmask = wmask; // @[Uncache.scala 96:24]
  assign io_out_req_bits_wen = wen; // @[Uncache.scala 86:24]
  assign io_out_req_bits_size = req_split ? 2'h2 : size; // @[Uncache.scala 97:30]
  assign io_out_resp_ready = state == 3'h2 | state == 3'h4; // @[Uncache.scala 89:47]
  always @(posedge clock) begin
    if (reset) begin // @[Uncache.scala 18:22]
      state <= 3'h0; // @[Uncache.scala 18:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        state <= 3'h1; // @[Uncache.scala 47:17]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Uncache.scala 52:29]
        state <= 3'h2; // @[Uncache.scala 53:15]
      end
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      state <= _GEN_11;
    end else begin
      state <= _GEN_19;
    end
    if (reset) begin // @[Uncache.scala 21:22]
      addr <= 32'h0; // @[Uncache.scala 21:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        addr <= io_in_req_bits_addr; // @[Uncache.scala 39:15]
      end
    end
    if (reset) begin // @[Uncache.scala 22:22]
      ren <= 1'h0; // @[Uncache.scala 22:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        ren <= io_in_req_bits_ren; // @[Uncache.scala 40:15]
      end
    end
    if (reset) begin // @[Uncache.scala 23:22]
      wdata <= 64'h0; // @[Uncache.scala 23:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        wdata <= io_in_req_bits_wdata; // @[Uncache.scala 41:15]
      end
    end
    if (reset) begin // @[Uncache.scala 24:22]
      wmask <= 8'h0; // @[Uncache.scala 24:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        wmask <= io_in_req_bits_wmask; // @[Uncache.scala 42:15]
      end
    end
    if (reset) begin // @[Uncache.scala 25:22]
      wen <= 1'h0; // @[Uncache.scala 25:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        wen <= io_in_req_bits_wen; // @[Uncache.scala 43:15]
      end
    end
    if (reset) begin // @[Uncache.scala 26:22]
      size <= 2'h0; // @[Uncache.scala 26:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        size <= io_in_req_bits_size; // @[Uncache.scala 44:15]
      end
    end
    if (reset) begin // @[Uncache.scala 29:24]
      rdata_1 <= 64'h0; // @[Uncache.scala 29:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        rdata_1 <= 64'h0; // @[Uncache.scala 45:17]
      end
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_4) begin // @[Conditional.scala 39:67]
        rdata_1 <= _GEN_10;
      end
    end
    if (reset) begin // @[Uncache.scala 30:24]
      rdata_2 <= 64'h0; // @[Uncache.scala 30:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Uncache.scala 38:28]
        rdata_2 <= 64'h0; // @[Uncache.scala 46:17]
      end
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        rdata_2 <= _GEN_20;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  ren = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  wdata = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  wmask = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  wen = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  size = _RAND_6[1:0];
  _RAND_7 = {2{`RANDOM}};
  rdata_1 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  rdata_2 = _RAND_8[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210340_CacheController_1(
  input         clock,
  input         reset, 
  output [5:0]   io_sram4_addr,
  output         io_sram4_cen,
  output         io_sram4_wen,
  output [127:0] io_sram4_wdata,
  input  [127:0] io_sram4_rdata,
  output [5:0]   io_sram5_addr,
  output         io_sram5_cen,
  output         io_sram5_wen,
  output [127:0] io_sram5_wdata,
  input  [127:0] io_sram5_rdata,
  output [5:0]   io_sram6_addr,
  output         io_sram6_cen,
  output         io_sram6_wen,
  output [127:0] io_sram6_wdata,
  input  [127:0] io_sram6_rdata,
  output [5:0]   io_sram7_addr,
  output         io_sram7_cen,
  output         io_sram7_wen,
  output [127:0] io_sram7_wdata,
  input  [127:0] io_sram7_rdata,    
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input         io_in_req_bits_ren,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input  [1:0]  io_in_req_bits_size,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_cache_req_ready,
  output        io_out_cache_req_valid,
  output [31:0] io_out_cache_req_bits_addr,
  output        io_out_cache_req_bits_aen,
  output        io_out_cache_req_bits_ren,
  output [63:0] io_out_cache_req_bits_wdata,
  output        io_out_cache_req_bits_wlast,
  output        io_out_cache_req_bits_wen,
  output        io_out_cache_resp_ready,
  input         io_out_cache_resp_valid,
  input  [63:0] io_out_cache_resp_bits_rdata,
  input         io_out_cache_resp_bits_rlast,
  input         io_out_uncache_req_ready,
  output        io_out_uncache_req_valid,
  output [31:0] io_out_uncache_req_bits_addr,
  output        io_out_uncache_req_bits_ren,
  output [63:0] io_out_uncache_req_bits_wdata,
  output [7:0]  io_out_uncache_req_bits_wmask,
  output        io_out_uncache_req_bits_wen,
  output [1:0]  io_out_uncache_req_bits_size,
  output        io_out_uncache_resp_ready,
  input         io_out_uncache_resp_valid,
  input  [63:0] io_out_uncache_resp_bits_rdata,
  input         fence_i,
  output        dcache_fi_complete
);

  wire [5:0] dcache_io_sram4_addr; 
  wire  dcache_io_sram4_cen; 
  wire  dcache_io_sram4_wen; 
  wire [127:0] dcache_io_sram4_wdata; 
  wire [127:0] dcache_io_sram4_rdata; 
  wire [5:0] dcache_io_sram5_addr; 
  wire  dcache_io_sram5_cen; 
  wire  dcache_io_sram5_wen; 
  wire [127:0] dcache_io_sram5_wdata; 
  wire [127:0] dcache_io_sram5_rdata; 
  wire [5:0] dcache_io_sram6_addr; 
  wire  dcache_io_sram6_cen; 
  wire  dcache_io_sram6_wen; 
  wire [127:0] dcache_io_sram6_wdata; 
  wire [127:0] dcache_io_sram6_rdata; 
  wire [5:0] dcache_io_sram7_addr; 
  wire  dcache_io_sram7_cen; 
  wire  dcache_io_sram7_wen; 
  wire [127:0] dcache_io_sram7_wdata; 
  wire [127:0] dcache_io_sram7_rdata;

  wire  cache_clock; // @[CacheController.scala 14:21]
  wire  cache_reset; // @[CacheController.scala 14:21]
  wire  cache_io_in_req_ready; // @[CacheController.scala 14:21]
  wire  cache_io_in_req_valid; // @[CacheController.scala 14:21]
  wire [31:0] cache_io_in_req_bits_addr; // @[CacheController.scala 14:21]
  wire [63:0] cache_io_in_req_bits_wdata; // @[CacheController.scala 14:21]
  wire [7:0] cache_io_in_req_bits_wmask; // @[CacheController.scala 14:21]
  wire  cache_io_in_req_bits_wen; // @[CacheController.scala 14:21]
  wire  cache_io_in_resp_ready; // @[CacheController.scala 14:21]
  wire  cache_io_in_resp_valid; // @[CacheController.scala 14:21]
  wire [63:0] cache_io_in_resp_bits_rdata; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_ready; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_valid; // @[CacheController.scala 14:21]
  wire [31:0] cache_io_out_req_bits_addr; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_bits_aen; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_bits_ren; // @[CacheController.scala 14:21]
  wire [63:0] cache_io_out_req_bits_wdata; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_bits_wlast; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_bits_wen; // @[CacheController.scala 14:21]
  wire  cache_io_out_resp_ready; // @[CacheController.scala 14:21]
  wire  cache_io_out_resp_valid; // @[CacheController.scala 14:21]
  wire [63:0] cache_io_out_resp_bits_rdata; // @[CacheController.scala 14:21]
  wire  cache_io_out_resp_bits_rlast; // @[CacheController.scala 14:21]
  wire  cache_fence_i_0; // @[CacheController.scala 14:21]
  wire  cache_dcache_fi_complete_0; // @[CacheController.scala 14:21]
  wire  uncache_clock; // @[CacheController.scala 15:23]
  wire  uncache_reset; // @[CacheController.scala 15:23]
  wire  uncache_io_in_req_ready; // @[CacheController.scala 15:23]
  wire  uncache_io_in_req_valid; // @[CacheController.scala 15:23]
  wire [31:0] uncache_io_in_req_bits_addr; // @[CacheController.scala 15:23]
  wire  uncache_io_in_req_bits_ren; // @[CacheController.scala 15:23]
  wire [63:0] uncache_io_in_req_bits_wdata; // @[CacheController.scala 15:23]
  wire [7:0] uncache_io_in_req_bits_wmask; // @[CacheController.scala 15:23]
  wire  uncache_io_in_req_bits_wen; // @[CacheController.scala 15:23]
  wire [1:0] uncache_io_in_req_bits_size; // @[CacheController.scala 15:23]
  wire  uncache_io_in_resp_ready; // @[CacheController.scala 15:23]
  wire  uncache_io_in_resp_valid; // @[CacheController.scala 15:23]
  wire [63:0] uncache_io_in_resp_bits_rdata; // @[CacheController.scala 15:23]
  wire  uncache_io_out_req_ready; // @[CacheController.scala 15:23]
  wire  uncache_io_out_req_valid; // @[CacheController.scala 15:23]
  wire [31:0] uncache_io_out_req_bits_addr; // @[CacheController.scala 15:23]
  wire  uncache_io_out_req_bits_ren; // @[CacheController.scala 15:23]
  wire [63:0] uncache_io_out_req_bits_wdata; // @[CacheController.scala 15:23]
  wire [7:0] uncache_io_out_req_bits_wmask; // @[CacheController.scala 15:23]
  wire  uncache_io_out_req_bits_wen; // @[CacheController.scala 15:23]
  wire [1:0] uncache_io_out_req_bits_size; // @[CacheController.scala 15:23]
  wire  uncache_io_out_resp_ready; // @[CacheController.scala 15:23]
  wire  uncache_io_out_resp_valid; // @[CacheController.scala 15:23]
  wire [63:0] uncache_io_out_resp_bits_rdata; // @[CacheController.scala 15:23]
  wire  crossbar1to2_clock; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_req_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_req_valid; // @[CacheController.scala 17:28]
  wire [31:0] crossbar1to2_io_in_req_bits_addr; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_req_bits_ren; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_in_req_bits_wdata; // @[CacheController.scala 17:28]
  wire [7:0] crossbar1to2_io_in_req_bits_wmask; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_req_bits_wen; // @[CacheController.scala 17:28]
  wire [1:0] crossbar1to2_io_in_req_bits_size; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_resp_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_resp_valid; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_in_resp_bits_rdata; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_req_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_req_valid; // @[CacheController.scala 17:28]
  wire [31:0] crossbar1to2_io_out_0_req_bits_addr; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_req_bits_ren; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_out_0_req_bits_wdata; // @[CacheController.scala 17:28]
  wire [7:0] crossbar1to2_io_out_0_req_bits_wmask; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_req_bits_wen; // @[CacheController.scala 17:28]
  wire [1:0] crossbar1to2_io_out_0_req_bits_size; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_resp_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_resp_valid; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_out_0_resp_bits_rdata; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_req_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_req_valid; // @[CacheController.scala 17:28]
  wire [31:0] crossbar1to2_io_out_1_req_bits_addr; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_req_bits_ren; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_out_1_req_bits_wdata; // @[CacheController.scala 17:28]
  wire [7:0] crossbar1to2_io_out_1_req_bits_wmask; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_req_bits_wen; // @[CacheController.scala 17:28]
  wire [1:0] crossbar1to2_io_out_1_req_bits_size; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_resp_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_resp_valid; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_out_1_resp_bits_rdata; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_to_1; // @[CacheController.scala 17:28]
  ysyx_210340_Cache_1 cache ( // @[CacheController.scala 14:21]
    .clock(cache_clock),
    .reset(cache_reset),
    .io_sram4_cen(dcache_io_sram4_cen), 
    .io_sram4_wen(dcache_io_sram4_wen), 
    .io_sram4_addr(dcache_io_sram4_addr), 
    .io_sram4_wdata(dcache_io_sram4_wdata), 
    .io_sram4_rdata(dcache_io_sram4_rdata), 
    .io_sram5_cen(dcache_io_sram5_cen), 
    .io_sram5_wen(dcache_io_sram5_wen), 
    .io_sram5_addr(dcache_io_sram5_addr), 
    .io_sram5_wdata(dcache_io_sram5_wdata), 
    .io_sram5_rdata(dcache_io_sram5_rdata), 
    .io_sram6_cen(dcache_io_sram6_cen), 
    .io_sram6_wen(dcache_io_sram6_wen), 
    .io_sram6_addr(dcache_io_sram6_addr), 
    .io_sram6_wdata(dcache_io_sram6_wdata), 
    .io_sram6_rdata(dcache_io_sram6_rdata),   
    .io_sram7_cen(dcache_io_sram7_cen), 
    .io_sram7_wen(dcache_io_sram7_wen), 
    .io_sram7_addr(dcache_io_sram7_addr), 
    .io_sram7_wdata(dcache_io_sram7_wdata), 
    .io_sram7_rdata(dcache_io_sram7_rdata),  
    .io_in_req_ready(cache_io_in_req_ready),
    .io_in_req_valid(cache_io_in_req_valid),
    .io_in_req_bits_addr(cache_io_in_req_bits_addr),
    .io_in_req_bits_wdata(cache_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(cache_io_in_req_bits_wmask),
    .io_in_req_bits_wen(cache_io_in_req_bits_wen),
    .io_in_resp_ready(cache_io_in_resp_ready),
    .io_in_resp_valid(cache_io_in_resp_valid),
    .io_in_resp_bits_rdata(cache_io_in_resp_bits_rdata),
    .io_out_req_ready(cache_io_out_req_ready),
    .io_out_req_valid(cache_io_out_req_valid),
    .io_out_req_bits_addr(cache_io_out_req_bits_addr),
    .io_out_req_bits_aen(cache_io_out_req_bits_aen),
    .io_out_req_bits_ren(cache_io_out_req_bits_ren),
    .io_out_req_bits_wdata(cache_io_out_req_bits_wdata),
    .io_out_req_bits_wlast(cache_io_out_req_bits_wlast),
    .io_out_req_bits_wen(cache_io_out_req_bits_wen),
    .io_out_resp_ready(cache_io_out_resp_ready),
    .io_out_resp_valid(cache_io_out_resp_valid),
    .io_out_resp_bits_rdata(cache_io_out_resp_bits_rdata),
    .io_out_resp_bits_rlast(cache_io_out_resp_bits_rlast),
    .fence_i_0(cache_fence_i_0),
    .dcache_fi_complete_0(cache_dcache_fi_complete_0)
  );

  assign io_sram4_addr = dcache_io_sram4_addr; // @[cpu.scala 167:22]
  assign io_sram4_cen = dcache_io_sram4_cen; // @[cpu.scala 167:22]
  assign io_sram4_wen = dcache_io_sram4_wen; // @[cpu.scala 167:22]
  assign io_sram4_wdata = dcache_io_sram4_wdata; // @[cpu.scala 167:22]
  assign io_sram5_addr = dcache_io_sram5_addr; // @[cpu.scala 168:22]
  assign io_sram5_cen = dcache_io_sram5_cen; // @[cpu.scala 168:22]
  assign io_sram5_wen = dcache_io_sram5_wen; // @[cpu.scala 168:22]
  assign io_sram5_wdata = dcache_io_sram5_wdata; // @[cpu.scala 168:22]
  assign io_sram6_addr = dcache_io_sram6_addr; // @[cpu.scala 169:22]
  assign io_sram6_cen = dcache_io_sram6_cen; // @[cpu.scala 169:22]
  assign io_sram6_wen = dcache_io_sram6_wen; // @[cpu.scala 169:22]
  assign io_sram6_wdata = dcache_io_sram6_wdata; // @[cpu.scala 169:22]
  assign io_sram7_addr = dcache_io_sram7_addr; // @[cpu.scala 170:22]
  assign io_sram7_cen = dcache_io_sram7_cen; // @[cpu.scala 170:22]
  assign io_sram7_wen = dcache_io_sram7_wen; // @[cpu.scala 170:22]
  assign io_sram7_wdata = dcache_io_sram7_wdata; // @[cpu.scala 170:22]

  assign dcache_io_sram4_rdata = io_sram4_rdata;
  assign dcache_io_sram5_rdata = io_sram5_rdata;
  assign dcache_io_sram6_rdata = io_sram6_rdata;
  assign dcache_io_sram7_rdata = io_sram7_rdata;

  ysyx_210340_Uncache_1 uncache ( // @[CacheController.scala 15:23]
    .clock(uncache_clock),
    .reset(uncache_reset),
    .io_in_req_ready(uncache_io_in_req_ready),
    .io_in_req_valid(uncache_io_in_req_valid),
    .io_in_req_bits_addr(uncache_io_in_req_bits_addr),
    .io_in_req_bits_ren(uncache_io_in_req_bits_ren),
    .io_in_req_bits_wdata(uncache_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(uncache_io_in_req_bits_wmask),
    .io_in_req_bits_wen(uncache_io_in_req_bits_wen),
    .io_in_req_bits_size(uncache_io_in_req_bits_size),
    .io_in_resp_ready(uncache_io_in_resp_ready),
    .io_in_resp_valid(uncache_io_in_resp_valid),
    .io_in_resp_bits_rdata(uncache_io_in_resp_bits_rdata),
    .io_out_req_ready(uncache_io_out_req_ready),
    .io_out_req_valid(uncache_io_out_req_valid),
    .io_out_req_bits_addr(uncache_io_out_req_bits_addr),
    .io_out_req_bits_ren(uncache_io_out_req_bits_ren),
    .io_out_req_bits_wdata(uncache_io_out_req_bits_wdata),
    .io_out_req_bits_wmask(uncache_io_out_req_bits_wmask),
    .io_out_req_bits_wen(uncache_io_out_req_bits_wen),
    .io_out_req_bits_size(uncache_io_out_req_bits_size),
    .io_out_resp_ready(uncache_io_out_resp_ready),
    .io_out_resp_valid(uncache_io_out_resp_valid),
    .io_out_resp_bits_rdata(uncache_io_out_resp_bits_rdata)
  );
  ysyx_210340_CacheBusCrossbar1to2 crossbar1to2 ( // @[CacheController.scala 17:28]
    .clock(crossbar1to2_clock),
    .io_in_req_ready(crossbar1to2_io_in_req_ready),
    .io_in_req_valid(crossbar1to2_io_in_req_valid),
    .io_in_req_bits_addr(crossbar1to2_io_in_req_bits_addr),
    .io_in_req_bits_ren(crossbar1to2_io_in_req_bits_ren),
    .io_in_req_bits_wdata(crossbar1to2_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(crossbar1to2_io_in_req_bits_wmask),
    .io_in_req_bits_wen(crossbar1to2_io_in_req_bits_wen),
    .io_in_req_bits_size(crossbar1to2_io_in_req_bits_size),
    .io_in_resp_ready(crossbar1to2_io_in_resp_ready),
    .io_in_resp_valid(crossbar1to2_io_in_resp_valid),
    .io_in_resp_bits_rdata(crossbar1to2_io_in_resp_bits_rdata),
    .io_out_0_req_ready(crossbar1to2_io_out_0_req_ready),
    .io_out_0_req_valid(crossbar1to2_io_out_0_req_valid),
    .io_out_0_req_bits_addr(crossbar1to2_io_out_0_req_bits_addr),
    .io_out_0_req_bits_ren(crossbar1to2_io_out_0_req_bits_ren),
    .io_out_0_req_bits_wdata(crossbar1to2_io_out_0_req_bits_wdata),
    .io_out_0_req_bits_wmask(crossbar1to2_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wen(crossbar1to2_io_out_0_req_bits_wen),
    .io_out_0_req_bits_size(crossbar1to2_io_out_0_req_bits_size),
    .io_out_0_resp_ready(crossbar1to2_io_out_0_resp_ready),
    .io_out_0_resp_valid(crossbar1to2_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(crossbar1to2_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(crossbar1to2_io_out_1_req_ready),
    .io_out_1_req_valid(crossbar1to2_io_out_1_req_valid),
    .io_out_1_req_bits_addr(crossbar1to2_io_out_1_req_bits_addr),
    .io_out_1_req_bits_ren(crossbar1to2_io_out_1_req_bits_ren),
    .io_out_1_req_bits_wdata(crossbar1to2_io_out_1_req_bits_wdata),
    .io_out_1_req_bits_wmask(crossbar1to2_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wen(crossbar1to2_io_out_1_req_bits_wen),
    .io_out_1_req_bits_size(crossbar1to2_io_out_1_req_bits_size),
    .io_out_1_resp_ready(crossbar1to2_io_out_1_resp_ready),
    .io_out_1_resp_valid(crossbar1to2_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(crossbar1to2_io_out_1_resp_bits_rdata),
    .io_to_1(crossbar1to2_io_to_1)
  );
  assign io_in_req_ready = crossbar1to2_io_in_req_ready; // @[CacheController.scala 19:22]
  assign io_in_resp_valid = crossbar1to2_io_in_resp_valid; // @[CacheController.scala 19:22]
  assign io_in_resp_bits_rdata = crossbar1to2_io_in_resp_bits_rdata; // @[CacheController.scala 19:22]
  assign io_out_cache_req_valid = cache_io_out_req_valid; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_addr = cache_io_out_req_bits_addr; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_aen = cache_io_out_req_bits_aen; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_ren = cache_io_out_req_bits_ren; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_wdata = cache_io_out_req_bits_wdata; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_wlast = cache_io_out_req_bits_wlast; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_wen = cache_io_out_req_bits_wen; // @[CacheController.scala 23:16]
  assign io_out_cache_resp_ready = cache_io_out_resp_ready; // @[CacheController.scala 23:16]
  assign io_out_uncache_req_valid = uncache_io_out_req_valid; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_addr = uncache_io_out_req_bits_addr; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_ren = uncache_io_out_req_bits_ren; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_wdata = uncache_io_out_req_bits_wdata; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_wmask = uncache_io_out_req_bits_wmask; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_wen = uncache_io_out_req_bits_wen; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_size = uncache_io_out_req_bits_size; // @[CacheController.scala 24:18]
  assign io_out_uncache_resp_ready = uncache_io_out_resp_ready; // @[CacheController.scala 24:18]
  assign dcache_fi_complete = cache_dcache_fi_complete_0;
  assign cache_clock = clock;
  assign cache_reset = reset;
  assign cache_io_in_req_valid = crossbar1to2_io_out_0_req_valid; // @[CacheController.scala 20:26]
  assign cache_io_in_req_bits_addr = crossbar1to2_io_out_0_req_bits_addr; // @[CacheController.scala 20:26]
  assign cache_io_in_req_bits_wdata = crossbar1to2_io_out_0_req_bits_wdata; // @[CacheController.scala 20:26]
  assign cache_io_in_req_bits_wmask = crossbar1to2_io_out_0_req_bits_wmask; // @[CacheController.scala 20:26]
  assign cache_io_in_req_bits_wen = crossbar1to2_io_out_0_req_bits_wen; // @[CacheController.scala 20:26]
  assign cache_io_in_resp_ready = crossbar1to2_io_out_0_resp_ready; // @[CacheController.scala 20:26]
  assign cache_io_out_req_ready = io_out_cache_req_ready; // @[CacheController.scala 23:16]
  assign cache_io_out_resp_valid = io_out_cache_resp_valid; // @[CacheController.scala 23:16]
  assign cache_io_out_resp_bits_rdata = io_out_cache_resp_bits_rdata; // @[CacheController.scala 23:16]
  assign cache_io_out_resp_bits_rlast = io_out_cache_resp_bits_rlast; // @[CacheController.scala 23:16]
  assign cache_fence_i_0 = fence_i;
  assign uncache_clock = clock;
  assign uncache_reset = reset;
  assign uncache_io_in_req_valid = crossbar1to2_io_out_1_req_valid; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_addr = crossbar1to2_io_out_1_req_bits_addr; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_ren = crossbar1to2_io_out_1_req_bits_ren; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_wdata = crossbar1to2_io_out_1_req_bits_wdata; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_wmask = crossbar1to2_io_out_1_req_bits_wmask; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_wen = crossbar1to2_io_out_1_req_bits_wen; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_size = crossbar1to2_io_out_1_req_bits_size; // @[CacheController.scala 21:26]
  assign uncache_io_in_resp_ready = crossbar1to2_io_out_1_resp_ready; // @[CacheController.scala 21:26]
  assign uncache_io_out_req_ready = io_out_uncache_req_ready; // @[CacheController.scala 24:18]
  assign uncache_io_out_resp_valid = io_out_uncache_resp_valid; // @[CacheController.scala 24:18]
  assign uncache_io_out_resp_bits_rdata = io_out_uncache_resp_bits_rdata; // @[CacheController.scala 24:18]
  assign crossbar1to2_clock = clock;
  assign crossbar1to2_io_in_req_valid = io_in_req_valid; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_addr = io_in_req_bits_addr; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_ren = io_in_req_bits_ren; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_wdata = io_in_req_bits_wdata; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_wmask = io_in_req_bits_wmask; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_wen = io_in_req_bits_wen; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_size = io_in_req_bits_size; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_resp_ready = io_in_resp_ready; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_out_0_req_ready = cache_io_in_req_ready; // @[CacheController.scala 20:26]
  assign crossbar1to2_io_out_0_resp_valid = cache_io_in_resp_valid; // @[CacheController.scala 20:26]
  assign crossbar1to2_io_out_0_resp_bits_rdata = cache_io_in_resp_bits_rdata; // @[CacheController.scala 20:26]
  assign crossbar1to2_io_out_1_req_ready = uncache_io_in_req_ready; // @[CacheController.scala 21:26]
  assign crossbar1to2_io_out_1_resp_valid = uncache_io_in_resp_valid; // @[CacheController.scala 21:26]
  assign crossbar1to2_io_out_1_resp_bits_rdata = uncache_io_in_resp_bits_rdata; // @[CacheController.scala 21:26]
  assign crossbar1to2_io_to_1 = ~io_in_req_bits_addr[31]; // @[CacheController.scala 13:45]
endmodule
module ysyx_210340_Clint(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input         io_in_req_bits_ren,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output        mtip_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtime; // @[Clint.scala 13:22]
  reg [63:0] mtimecmp; // @[Clint.scala 14:25]
  wire [63:0] _mtime_T_1 = mtime + 64'ha; // @[Clint.scala 24:18]
  wire [15:0] clint_addr = io_in_req_bits_addr[15:0]; // @[Clint.scala 26:39]
  wire  _clint_ren_T = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  wire  clint_ren = io_in_req_bits_ren & _clint_ren_T; // @[Clint.scala 28:38]
  wire [7:0] clint_wmask_lo_lo_lo = io_in_req_bits_wmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] clint_wmask_lo_lo_hi = io_in_req_bits_wmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] clint_wmask_lo_hi_lo = io_in_req_bits_wmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] clint_wmask_lo_hi_hi = io_in_req_bits_wmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] clint_wmask_hi_lo_lo = io_in_req_bits_wmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] clint_wmask_hi_lo_hi = io_in_req_bits_wmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] clint_wmask_hi_hi_lo = io_in_req_bits_wmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] clint_wmask_hi_hi_hi = io_in_req_bits_wmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] clint_wmask = {clint_wmask_hi_hi_hi,clint_wmask_hi_hi_lo,clint_wmask_hi_lo_hi,clint_wmask_hi_lo_lo,
    clint_wmask_lo_hi_hi,clint_wmask_lo_hi_lo,clint_wmask_lo_lo_hi,clint_wmask_lo_lo_lo}; // @[Cat.scala 30:58]
  wire  clint_wen = io_in_req_bits_wen & _clint_ren_T; // @[Clint.scala 31:38]
  wire  _T_1 = clint_addr == 16'h4000; // @[Clint.scala 33:26]
  wire  _T_4 = clint_addr == 16'hbff8; // @[Clint.scala 35:33]
  wire [63:0] _GEN_0 = clint_addr == 16'hbff8 & clint_ren ? mtime : 64'h0; // @[Clint.scala 35:61 Clint.scala 36:17 Clint.scala 38:17]
  wire [63:0] _mtimecmp_T = io_in_req_bits_wdata & clint_wmask; // @[Clint.scala 42:30]
  reg [63:0] reg_rdata; // @[Clint.scala 47:26]
  reg [1:0] state; // @[Clint.scala 49:22]
  wire  _T_12 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_13 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_14 = io_in_resp_ready & io_in_resp_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_8 = _T_14 ? 2'h0 : state; // @[Clint.scala 61:32 Clint.scala 62:15 Clint.scala 49:22]
  wire  _T_15 = 2'h2 == state; // @[Conditional.scala 37:30]
  reg  mtip; // @[Clint.scala 79:21]
  assign io_in_req_ready = state == 2'h0; // @[Clint.scala 72:29]
  assign io_in_resp_valid = state != 2'h0; // @[Clint.scala 73:30]
  assign io_in_resp_bits_rdata = reg_rdata; // @[Clint.scala 75:25]
  assign mtip_0 = mtip;
  always @(posedge clock) begin
    if (reset) begin // @[Clint.scala 13:22]
      mtime <= 64'h0; // @[Clint.scala 13:22]
    end else if (_T_1 & clint_wen) begin // @[Clint.scala 41:54]
      mtime <= _mtime_T_1; // @[Clint.scala 24:9]
    end else if (_T_4 & clint_wen) begin // @[Clint.scala 43:61]
      mtime <= _mtimecmp_T; // @[Clint.scala 44:11]
    end else begin
      mtime <= _mtime_T_1; // @[Clint.scala 24:9]
    end
    if (reset) begin // @[Clint.scala 14:25]
      mtimecmp <= 64'h0; // @[Clint.scala 14:25]
    end else if (_T_1 & clint_wen) begin // @[Clint.scala 41:54]
      mtimecmp <= _mtimecmp_T; // @[Clint.scala 42:14]
    end
    if (reset) begin // @[Clint.scala 47:26]
      reg_rdata <= 64'h0; // @[Clint.scala 47:26]
    end else if (_T_12) begin // @[Conditional.scala 40:58]
      if (clint_ren) begin // @[Clint.scala 53:24]
        if (clint_addr == 16'h4000 & clint_ren) begin // @[Clint.scala 33:54]
          reg_rdata <= mtimecmp; // @[Clint.scala 34:17]
        end else begin
          reg_rdata <= _GEN_0;
        end
      end
    end
    if (reset) begin // @[Clint.scala 49:22]
      state <= 2'h0; // @[Clint.scala 49:22]
    end else if (_T_12) begin // @[Conditional.scala 40:58]
      if (clint_ren) begin // @[Clint.scala 53:24]
        state <= 2'h1; // @[Clint.scala 55:15]
      end else if (clint_wen) begin // @[Clint.scala 56:31]
        state <= 2'h2; // @[Clint.scala 57:15]
      end
    end else if (_T_13) begin // @[Conditional.scala 39:67]
      state <= _GEN_8;
    end else if (_T_15) begin // @[Conditional.scala 39:67]
      state <= _GEN_8;
    end
    if (reset) begin // @[Clint.scala 79:21]
      mtip <= 1'h0; // @[Clint.scala 79:21]
    end else begin
      mtip <= mtime >= mtimecmp; // @[Clint.scala 80:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtime = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtimecmp = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  reg_rdata = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  mtip = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210340_Core(
  input         clock,
  input         reset,
  output [5:0]   io_sram0_addr,
  output         io_sram0_cen,
  output         io_sram0_wen,
  output [127:0] io_sram0_wdata,
  input  [127:0] io_sram0_rdata,
  output [5:0]   io_sram1_addr,
  output         io_sram1_cen,
  output         io_sram1_wen,
  output [127:0] io_sram1_wdata,
  input  [127:0] io_sram1_rdata,
  output [5:0]   io_sram2_addr,
  output         io_sram2_cen,
  output         io_sram2_wen,
  output [127:0] io_sram2_wdata,
  input  [127:0] io_sram2_rdata,
  output [5:0]   io_sram3_addr,
  output         io_sram3_cen,
  output         io_sram3_wen,
  output [127:0] io_sram3_wdata,
  input  [127:0] io_sram3_rdata,
  output [5:0]   io_sram4_addr,
  output         io_sram4_cen,
  output         io_sram4_wen,
  output [127:0] io_sram4_wdata,
  input  [127:0] io_sram4_rdata,
  output [5:0]   io_sram5_addr,
  output         io_sram5_cen,
  output         io_sram5_wen,
  output [127:0] io_sram5_wdata,
  input  [127:0] io_sram5_rdata,
  output [5:0]   io_sram6_addr,
  output         io_sram6_cen,
  output         io_sram6_wen,
  output [127:0] io_sram6_wdata,
  input  [127:0] io_sram6_rdata,
  output [5:0]   io_sram7_addr,
  output         io_sram7_cen,
  output         io_sram7_wen,
  output [127:0] io_sram7_wdata,
  input  [127:0] io_sram7_rdata,  
  input         io_core_bus_0_req_ready,
  output        io_core_bus_0_req_valid,
  output [31:0] io_core_bus_0_req_bits_addr,
  output        io_core_bus_0_req_bits_aen,
  output        io_core_bus_0_req_bits_ren,
  output [63:0] io_core_bus_0_req_bits_wdata,
  output        io_core_bus_0_req_bits_wlast,
  output        io_core_bus_0_req_bits_wen,
  output        io_core_bus_0_resp_ready,
  input         io_core_bus_0_resp_valid,
  input  [63:0] io_core_bus_0_resp_bits_rdata,
  input         io_core_bus_0_resp_bits_rlast,
  input         io_core_bus_1_req_ready,
  output        io_core_bus_1_req_valid,
  output [31:0] io_core_bus_1_req_bits_addr,
  output        io_core_bus_1_req_bits_aen,
  output        io_core_bus_1_req_bits_ren,
  output [63:0] io_core_bus_1_req_bits_wdata,
  output        io_core_bus_1_req_bits_wlast,
  output        io_core_bus_1_req_bits_wen,
  output        io_core_bus_1_resp_ready,
  input         io_core_bus_1_resp_valid,
  input  [63:0] io_core_bus_1_resp_bits_rdata,
  input         io_core_bus_1_resp_bits_rlast,
  input         io_core_bus_2_req_ready,
  output        io_core_bus_2_req_valid,
  output [31:0] io_core_bus_2_req_bits_addr,
  output        io_core_bus_2_req_bits_ren,
  output [63:0] io_core_bus_2_req_bits_wdata,
  output [7:0]  io_core_bus_2_req_bits_wmask,
  output        io_core_bus_2_req_bits_wen,
  output [1:0]  io_core_bus_2_req_bits_size,
  output        io_core_bus_2_resp_ready,
  input         io_core_bus_2_resp_valid,
  input  [63:0] io_core_bus_2_resp_bits_rdata,
  input         io_core_bus_3_req_ready,
  output        io_core_bus_3_req_valid,
  output [31:0] io_core_bus_3_req_bits_addr,
  output        io_core_bus_3_req_bits_ren,
  output [63:0] io_core_bus_3_req_bits_wdata,
  output [7:0]  io_core_bus_3_req_bits_wmask,
  output        io_core_bus_3_req_bits_wen,
  output [1:0]  io_core_bus_3_req_bits_size,
  output        io_core_bus_3_resp_ready,
  input         io_core_bus_3_resp_valid,
  input  [63:0] io_core_bus_3_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  fetch_clock; // @[Core.scala 18:21]
  wire  fetch_reset; // @[Core.scala 18:21]
  wire  fetch_io_stall; // @[Core.scala 18:21]
  wire  fetch_io_flush; // @[Core.scala 18:21]
  wire  fetch_io_br_en; // @[Core.scala 18:21]
  wire [31:0] fetch_io_br_addr; // @[Core.scala 18:21]
  wire [31:0] fetch_io_out_pc; // @[Core.scala 18:21]
  wire [31:0] fetch_io_out_inst; // @[Core.scala 18:21]
  wire  fetch_io_out_imem_hs; // @[Core.scala 18:21]
  wire  fetch_io_imem_req_ready; // @[Core.scala 18:21]
  wire  fetch_io_imem_req_valid; // @[Core.scala 18:21]
  wire [31:0] fetch_io_imem_req_bits_addr; // @[Core.scala 18:21]
  wire  fetch_io_imem_resp_ready; // @[Core.scala 18:21]
  wire  fetch_io_imem_resp_valid; // @[Core.scala 18:21]
  wire [63:0] fetch_io_imem_resp_bits_rdata; // @[Core.scala 18:21]
  wire  icache_clock; // @[Core.scala 20:22]
  wire  icache_reset; // @[Core.scala 20:22]
  wire  icache_io_in_req_ready; // @[Core.scala 20:22]
  wire  icache_io_in_req_valid; // @[Core.scala 20:22]
  wire [31:0] icache_io_in_req_bits_addr; // @[Core.scala 20:22]
  wire  icache_io_in_resp_ready; // @[Core.scala 20:22]
  wire  icache_io_in_resp_valid; // @[Core.scala 20:22]
  wire [63:0] icache_io_in_resp_bits_rdata; // @[Core.scala 20:22]
  wire  icache_io_out_cache_req_ready; // @[Core.scala 20:22]
  wire  icache_io_out_cache_req_valid; // @[Core.scala 20:22]
  wire [31:0] icache_io_out_cache_req_bits_addr; // @[Core.scala 20:22]
  wire  icache_io_out_cache_req_bits_aen; // @[Core.scala 20:22]
  wire  icache_io_out_cache_req_bits_ren; // @[Core.scala 20:22]
  wire [63:0] icache_io_out_cache_req_bits_wdata; // @[Core.scala 20:22]
  wire  icache_io_out_cache_req_bits_wlast; // @[Core.scala 20:22]
  wire  icache_io_out_cache_req_bits_wen; // @[Core.scala 20:22]
  wire  icache_io_out_cache_resp_ready; // @[Core.scala 20:22]
  wire  icache_io_out_cache_resp_valid; // @[Core.scala 20:22]
  wire [63:0] icache_io_out_cache_resp_bits_rdata; // @[Core.scala 20:22]
  wire  icache_io_out_cache_resp_bits_rlast; // @[Core.scala 20:22]
  wire  icache_io_out_uncache_req_ready; // @[Core.scala 20:22]
  wire  icache_io_out_uncache_req_valid; // @[Core.scala 20:22]
  wire [31:0] icache_io_out_uncache_req_bits_addr; // @[Core.scala 20:22]
  wire  icache_io_out_uncache_req_bits_ren; // @[Core.scala 20:22]
  wire [63:0] icache_io_out_uncache_req_bits_wdata; // @[Core.scala 20:22]
  wire [7:0] icache_io_out_uncache_req_bits_wmask; // @[Core.scala 20:22]
  wire  icache_io_out_uncache_req_bits_wen; // @[Core.scala 20:22]
  wire [1:0] icache_io_out_uncache_req_bits_size; // @[Core.scala 20:22]
  wire  icache_io_out_uncache_resp_ready; // @[Core.scala 20:22]
  wire  icache_io_out_uncache_resp_valid; // @[Core.scala 20:22]
  wire [63:0] icache_io_out_uncache_resp_bits_rdata; // @[Core.scala 20:22]
  wire  icache_fence_i; // @[Core.scala 20:22]
  wire  icache_dcache_fi_complete; // @[Core.scala 20:22]
  wire  if_id_reg_clock; // @[Core.scala 25:25]
  wire  if_id_reg_reset; // @[Core.scala 25:25]
  wire [31:0] if_id_reg_io_in_pc; // @[Core.scala 25:25]
  wire [31:0] if_id_reg_io_in_inst; // @[Core.scala 25:25]
  wire  if_id_reg_io_in_imem_hs; // @[Core.scala 25:25]
  wire [31:0] if_id_reg_io_out_pc; // @[Core.scala 25:25]
  wire [31:0] if_id_reg_io_out_inst; // @[Core.scala 25:25]
  wire  if_id_reg_io_out_imem_hs; // @[Core.scala 25:25]
  wire  if_id_reg_io_flush; // @[Core.scala 25:25]
  wire  if_id_reg_io_stall; // @[Core.scala 25:25]
  wire [31:0] decode_io_inst; // @[Core.scala 30:22]
  wire [4:0] decode_io_rs1_addr; // @[Core.scala 30:22]
  wire [1:0] decode_io_rs1_type; // @[Core.scala 30:22]
  wire [4:0] decode_io_rs2_addr; // @[Core.scala 30:22]
  wire [1:0] decode_io_rs2_type; // @[Core.scala 30:22]
  wire [4:0] decode_io_rd_addr; // @[Core.scala 30:22]
  wire  decode_io_rd_en; // @[Core.scala 30:22]
  wire [5:0] decode_io_op_type; // @[Core.scala 30:22]
  wire [2:0] decode_io_fuType; // @[Core.scala 30:22]
  wire [63:0] decode_io_imm; // @[Core.scala 30:22]
  wire [63:0] decode_io_csr_imm; // @[Core.scala 30:22]
  wire  rf_clock; // @[Core.scala 33:18]
  wire  rf_reset; // @[Core.scala 33:18]
  wire [31:0] rf_io_pc; // @[Core.scala 33:18]
  wire [4:0] rf_io_rs1_addr; // @[Core.scala 33:18]
  wire [4:0] rf_io_rs2_addr; // @[Core.scala 33:18]
  wire [1:0] rf_io_rs1_type; // @[Core.scala 33:18]
  wire [1:0] rf_io_rs2_type; // @[Core.scala 33:18]
  wire [4:0] rf_io_rd_addr; // @[Core.scala 33:18]
  wire  rf_io_rd_en; // @[Core.scala 33:18]
  wire [63:0] rf_io_rd_data; // @[Core.scala 33:18]
  wire [63:0] rf_io_imm; // @[Core.scala 33:18]
  wire [63:0] rf_io_csr_imm; // @[Core.scala 33:18]
  wire  rf_io_irq; // @[Core.scala 33:18]
  wire [63:0] rf_io_rs1; // @[Core.scala 33:18]
  wire [63:0] rf_io_rs2; // @[Core.scala 33:18]
  wire [63:0] rf_io_src2; // @[Core.scala 33:18]
  wire [31:0] execution_io_pc; // @[Core.scala 42:25]
  wire [5:0] execution_io_op_type; // @[Core.scala 42:25]
  wire [63:0] execution_io_rs1; // @[Core.scala 42:25]
  wire [63:0] execution_io_rs2; // @[Core.scala 42:25]
  wire [63:0] execution_io_src2; // @[Core.scala 42:25]
  wire [2:0] execution_io_fuType; // @[Core.scala 42:25]
  wire [63:0] execution_io_imm; // @[Core.scala 42:25]
  wire [31:0] execution_io_csr_Jmp_addr; // @[Core.scala 42:25]
  wire  execution_io_csr_Jmp_en; // @[Core.scala 42:25]
  wire [63:0] execution_io_csr_data; // @[Core.scala 42:25]
  wire  execution_io_br_en; // @[Core.scala 42:25]
  wire [31:0] execution_io_br_addr; // @[Core.scala 42:25]
  wire [63:0] execution_io_rd_data; // @[Core.scala 42:25]
  wire  execution_fence_i_0; // @[Core.scala 42:25]
  wire  id_ex_reg_clock; // @[Core.scala 49:25]
  wire  id_ex_reg_reset; // @[Core.scala 49:25]
  wire [31:0] id_ex_reg_io_in_pc; // @[Core.scala 49:25]
  wire  id_ex_reg_io_in_br_en; // @[Core.scala 49:25]
  wire [31:0] id_ex_reg_io_in_br_addr; // @[Core.scala 49:25]
  wire [5:0] id_ex_reg_io_in_op_type; // @[Core.scala 49:25]
  wire [2:0] id_ex_reg_io_in_fuType; // @[Core.scala 49:25]
  wire [63:0] id_ex_reg_io_in_rs1; // @[Core.scala 49:25]
  wire [63:0] id_ex_reg_io_in_rs2; // @[Core.scala 49:25]
  wire [4:0] id_ex_reg_io_in_rd_addr; // @[Core.scala 49:25]
  wire [63:0] id_ex_reg_io_in_src2; // @[Core.scala 49:25]
  wire  id_ex_reg_io_in_rd_en; // @[Core.scala 49:25]
  wire  id_ex_reg_io_in_imem_hs; // @[Core.scala 49:25]
  wire [63:0] id_ex_reg_io_in_rd_data; // @[Core.scala 49:25]
  wire [31:0] id_ex_reg_io_out_pc; // @[Core.scala 49:25]
  wire  id_ex_reg_io_out_br_en; // @[Core.scala 49:25]
  wire [31:0] id_ex_reg_io_out_br_addr; // @[Core.scala 49:25]
  wire [5:0] id_ex_reg_io_out_op_type; // @[Core.scala 49:25]
  wire [2:0] id_ex_reg_io_out_fuType; // @[Core.scala 49:25]
  wire [63:0] id_ex_reg_io_out_rs1; // @[Core.scala 49:25]
  wire [63:0] id_ex_reg_io_out_rs2; // @[Core.scala 49:25]
  wire [4:0] id_ex_reg_io_out_rd_addr; // @[Core.scala 49:25]
  wire [63:0] id_ex_reg_io_out_src2; // @[Core.scala 49:25]
  wire  id_ex_reg_io_out_rd_en; // @[Core.scala 49:25]
  wire  id_ex_reg_io_out_imem_hs; // @[Core.scala 49:25]
  wire [63:0] id_ex_reg_io_out_rd_data; // @[Core.scala 49:25]
  wire  id_ex_reg_io_stall; // @[Core.scala 49:25]
  wire  mem_clock; // @[Core.scala 67:19]
  wire  mem_reset; // @[Core.scala 67:19]
  wire [31:0] mem_io_pc; // @[Core.scala 67:19]
  wire [5:0] mem_io_op_type; // @[Core.scala 67:19]
  wire [63:0] mem_io_rs1; // @[Core.scala 67:19]
  wire [63:0] mem_io_rs2; // @[Core.scala 67:19]
  wire [63:0] mem_io_src2; // @[Core.scala 67:19]
  wire [2:0] mem_io_fuType; // @[Core.scala 67:19]
  wire  mem_io_irq; // @[Core.scala 67:19]
  wire  mem_io_mem_en; // @[Core.scala 67:19]
  wire [63:0] mem_io_rd_data; // @[Core.scala 67:19]
  wire  mem_io_busy; // @[Core.scala 67:19]
  wire  mem_io_dmem_hs; // @[Core.scala 67:19]
  wire  mem_io_resp_success; // @[Core.scala 67:19]
  wire  mem_io_dmem_req_ready; // @[Core.scala 67:19]
  wire  mem_io_dmem_req_valid; // @[Core.scala 67:19]
  wire [31:0] mem_io_dmem_req_bits_addr; // @[Core.scala 67:19]
  wire  mem_io_dmem_req_bits_ren; // @[Core.scala 67:19]
  wire [63:0] mem_io_dmem_req_bits_wdata; // @[Core.scala 67:19]
  wire [7:0] mem_io_dmem_req_bits_wmask; // @[Core.scala 67:19]
  wire  mem_io_dmem_req_bits_wen; // @[Core.scala 67:19]
  wire [1:0] mem_io_dmem_req_bits_size; // @[Core.scala 67:19]
  wire  mem_io_dmem_resp_ready; // @[Core.scala 67:19]
  wire  mem_io_dmem_resp_valid; // @[Core.scala 67:19]
  wire [63:0] mem_io_dmem_resp_bits_rdata; // @[Core.scala 67:19]
  wire  csr_clock; // @[Core.scala 77:19]
  wire  csr_reset; // @[Core.scala 77:19]
  wire [31:0] csr_io_pc; // @[Core.scala 77:19]
  wire [2:0] csr_io_fuType; // @[Core.scala 77:19]
  wire [5:0] csr_io_op_type; // @[Core.scala 77:19]
  wire [63:0] csr_io_rs1; // @[Core.scala 77:19]
  wire [63:0] csr_io_rs2; // @[Core.scala 77:19]
  wire  csr_io_if_valid; // @[Core.scala 77:19]
  wire  csr_io_mem_en; // @[Core.scala 77:19]
  wire  csr_io_mem_valid; // @[Core.scala 77:19]
  wire [31:0] csr_io_csr_Jmp_addr; // @[Core.scala 77:19]
  wire  csr_io_csr_Jmp_en; // @[Core.scala 77:19]
  wire [63:0] csr_io_csr_data; // @[Core.scala 77:19]
  wire  csr_io_irq; // @[Core.scala 77:19]
  wire  csr_mtip_0; // @[Core.scala 77:19]
  wire  crossbar1to2_clock; // @[Core.scala 87:28]
  wire  crossbar1to2_io_in_req_ready; // @[Core.scala 87:28]
  wire  crossbar1to2_io_in_req_valid; // @[Core.scala 87:28]
  wire [31:0] crossbar1to2_io_in_req_bits_addr; // @[Core.scala 87:28]
  wire  crossbar1to2_io_in_req_bits_ren; // @[Core.scala 87:28]
  wire [63:0] crossbar1to2_io_in_req_bits_wdata; // @[Core.scala 87:28]
  wire [7:0] crossbar1to2_io_in_req_bits_wmask; // @[Core.scala 87:28]
  wire  crossbar1to2_io_in_req_bits_wen; // @[Core.scala 87:28]
  wire [1:0] crossbar1to2_io_in_req_bits_size; // @[Core.scala 87:28]
  wire  crossbar1to2_io_in_resp_ready; // @[Core.scala 87:28]
  wire  crossbar1to2_io_in_resp_valid; // @[Core.scala 87:28]
  wire [63:0] crossbar1to2_io_in_resp_bits_rdata; // @[Core.scala 87:28]
  wire  crossbar1to2_io_out_0_req_ready; // @[Core.scala 87:28]
  wire  crossbar1to2_io_out_0_req_valid; // @[Core.scala 87:28]
  wire [31:0] crossbar1to2_io_out_0_req_bits_addr; // @[Core.scala 87:28]
  wire  crossbar1to2_io_out_0_req_bits_ren; // @[Core.scala 87:28]
  wire [63:0] crossbar1to2_io_out_0_req_bits_wdata; // @[Core.scala 87:28]
  wire [7:0] crossbar1to2_io_out_0_req_bits_wmask; // @[Core.scala 87:28]
  wire  crossbar1to2_io_out_0_req_bits_wen; // @[Core.scala 87:28]
  wire [1:0] crossbar1to2_io_out_0_req_bits_size; // @[Core.scala 87:28]
  wire  crossbar1to2_io_out_0_resp_ready; // @[Core.scala 87:28]
  wire  crossbar1to2_io_out_0_resp_valid; // @[Core.scala 87:28]
  wire [63:0] crossbar1to2_io_out_0_resp_bits_rdata; // @[Core.scala 87:28]
  wire  crossbar1to2_io_out_1_req_ready; // @[Core.scala 87:28]
  wire  crossbar1to2_io_out_1_req_valid; // @[Core.scala 87:28]
  wire [31:0] crossbar1to2_io_out_1_req_bits_addr; // @[Core.scala 87:28]
  wire  crossbar1to2_io_out_1_req_bits_ren; // @[Core.scala 87:28]
  wire [63:0] crossbar1to2_io_out_1_req_bits_wdata; // @[Core.scala 87:28]
  wire [7:0] crossbar1to2_io_out_1_req_bits_wmask; // @[Core.scala 87:28]
  wire  crossbar1to2_io_out_1_req_bits_wen; // @[Core.scala 87:28]
  wire [1:0] crossbar1to2_io_out_1_req_bits_size; // @[Core.scala 87:28]
  wire  crossbar1to2_io_out_1_resp_ready; // @[Core.scala 87:28]
  wire  crossbar1to2_io_out_1_resp_valid; // @[Core.scala 87:28]
  wire [63:0] crossbar1to2_io_out_1_resp_bits_rdata; // @[Core.scala 87:28]
  wire  crossbar1to2_io_to_1; // @[Core.scala 87:28]
  wire  dcache_clock; // @[Core.scala 94:22]
  wire  dcache_reset; // @[Core.scala 94:22]
  wire  dcache_io_in_req_ready; // @[Core.scala 94:22]
  wire  dcache_io_in_req_valid; // @[Core.scala 94:22]
  wire [31:0] dcache_io_in_req_bits_addr; // @[Core.scala 94:22]
  wire  dcache_io_in_req_bits_ren; // @[Core.scala 94:22]
  wire [63:0] dcache_io_in_req_bits_wdata; // @[Core.scala 94:22]
  wire [7:0] dcache_io_in_req_bits_wmask; // @[Core.scala 94:22]
  wire  dcache_io_in_req_bits_wen; // @[Core.scala 94:22]
  wire [1:0] dcache_io_in_req_bits_size; // @[Core.scala 94:22]
  wire  dcache_io_in_resp_ready; // @[Core.scala 94:22]
  wire  dcache_io_in_resp_valid; // @[Core.scala 94:22]
  wire [63:0] dcache_io_in_resp_bits_rdata; // @[Core.scala 94:22]
  wire  dcache_io_out_cache_req_ready; // @[Core.scala 94:22]
  wire  dcache_io_out_cache_req_valid; // @[Core.scala 94:22]
  wire [31:0] dcache_io_out_cache_req_bits_addr; // @[Core.scala 94:22]
  wire  dcache_io_out_cache_req_bits_aen; // @[Core.scala 94:22]
  wire  dcache_io_out_cache_req_bits_ren; // @[Core.scala 94:22]
  wire [63:0] dcache_io_out_cache_req_bits_wdata; // @[Core.scala 94:22]
  wire  dcache_io_out_cache_req_bits_wlast; // @[Core.scala 94:22]
  wire  dcache_io_out_cache_req_bits_wen; // @[Core.scala 94:22]
  wire  dcache_io_out_cache_resp_ready; // @[Core.scala 94:22]
  wire  dcache_io_out_cache_resp_valid; // @[Core.scala 94:22]
  wire [63:0] dcache_io_out_cache_resp_bits_rdata; // @[Core.scala 94:22]
  wire  dcache_io_out_cache_resp_bits_rlast; // @[Core.scala 94:22]
  wire  dcache_io_out_uncache_req_ready; // @[Core.scala 94:22]
  wire  dcache_io_out_uncache_req_valid; // @[Core.scala 94:22]
  wire [31:0] dcache_io_out_uncache_req_bits_addr; // @[Core.scala 94:22]
  wire  dcache_io_out_uncache_req_bits_ren; // @[Core.scala 94:22]
  wire [63:0] dcache_io_out_uncache_req_bits_wdata; // @[Core.scala 94:22]
  wire [7:0] dcache_io_out_uncache_req_bits_wmask; // @[Core.scala 94:22]
  wire  dcache_io_out_uncache_req_bits_wen; // @[Core.scala 94:22]
  wire [1:0] dcache_io_out_uncache_req_bits_size; // @[Core.scala 94:22]
  wire  dcache_io_out_uncache_resp_ready; // @[Core.scala 94:22]
  wire  dcache_io_out_uncache_resp_valid; // @[Core.scala 94:22]
  wire [63:0] dcache_io_out_uncache_resp_bits_rdata; // @[Core.scala 94:22]
  wire  dcache_fence_i; // @[Core.scala 94:22]
  wire  dcache_dcache_fi_complete; // @[Core.scala 94:22]
  wire  clint_clock; // @[Core.scala 99:21]
  wire  clint_reset; // @[Core.scala 99:21]
  wire  clint_io_in_req_ready; // @[Core.scala 99:21]
  wire  clint_io_in_req_valid; // @[Core.scala 99:21]
  wire [31:0] clint_io_in_req_bits_addr; // @[Core.scala 99:21]
  wire  clint_io_in_req_bits_ren; // @[Core.scala 99:21]
  wire [63:0] clint_io_in_req_bits_wdata; // @[Core.scala 99:21]
  wire [7:0] clint_io_in_req_bits_wmask; // @[Core.scala 99:21]
  wire  clint_io_in_req_bits_wen; // @[Core.scala 99:21]
  wire  clint_io_in_resp_ready; // @[Core.scala 99:21]
  wire  clint_io_in_resp_valid; // @[Core.scala 99:21]
  wire [63:0] clint_io_in_resp_bits_rdata; // @[Core.scala 99:21]
  wire  clint_mtip_0; // @[Core.scala 99:21]
  wire  _reg_wen_T_2 = mem_io_mem_en & ~id_ex_reg_io_out_op_type[3]; // @[Core.scala 75:35]
  reg  reg_wen_REG; // @[Core.scala 75:85]
  wire [63:0] _rf_io_rd_data_T_4 = _reg_wen_T_2 ? mem_io_rd_data : id_ex_reg_io_out_rd_data; // @[Core.scala 108:87]

  wire [5:0] icache_io_sram0_addr; 
  wire  icache_io_sram0_cen; 
  wire  icache_io_sram0_wen; 
  wire [127:0] icache_io_sram0_wdata; 
  wire [127:0] icache_io_sram0_rdata; 
  wire [5:0] icache_io_sram1_addr; 
  wire  icache_io_sram1_cen; 
  wire  icache_io_sram1_wen; 
  wire [127:0] icache_io_sram1_wdata; 
  wire [127:0] icache_io_sram1_rdata; 
  wire [5:0] icache_io_sram2_addr; 
  wire  icache_io_sram2_cen; 
  wire  icache_io_sram2_wen; 
  wire [127:0] icache_io_sram2_wdata; 
  wire [127:0] icache_io_sram2_rdata; 
  wire [5:0] icache_io_sram3_addr; 
  wire  icache_io_sram3_cen; 
  wire  icache_io_sram3_wen; 
  wire [127:0] icache_io_sram3_wdata; 
  wire [127:0] icache_io_sram3_rdata; 
  wire [5:0] dcache_io_sram4_addr; 
  wire  dcache_io_sram4_cen; 
  wire  dcache_io_sram4_wen; 
  wire [127:0] dcache_io_sram4_wdata; 
  wire [127:0] dcache_io_sram4_rdata; 
  wire [5:0] dcache_io_sram5_addr; 
  wire  dcache_io_sram5_cen; 
  wire  dcache_io_sram5_wen; 
  wire [127:0] dcache_io_sram5_wdata; 
  wire [127:0] dcache_io_sram5_rdata; 
  wire [5:0] dcache_io_sram6_addr; 
  wire  dcache_io_sram6_cen; 
  wire  dcache_io_sram6_wen; 
  wire [127:0] dcache_io_sram6_wdata; 
  wire [127:0] dcache_io_sram6_rdata; 
  wire [5:0] dcache_io_sram7_addr; 
  wire  dcache_io_sram7_cen; 
  wire  dcache_io_sram7_wen; 
  wire [127:0] dcache_io_sram7_wdata; 
  wire [127:0] dcache_io_sram7_rdata; 

  ysyx_210340_InstFetch fetch ( // @[Core.scala 18:21]
    .clock(fetch_clock),
    .reset(fetch_reset),
    .io_stall(fetch_io_stall),
    .io_flush(fetch_io_flush),
    .io_br_en(fetch_io_br_en),
    .io_br_addr(fetch_io_br_addr),
    .io_out_pc(fetch_io_out_pc),
    .io_out_inst(fetch_io_out_inst),
    .io_out_imem_hs(fetch_io_out_imem_hs),
    .io_imem_req_ready(fetch_io_imem_req_ready),
    .io_imem_req_valid(fetch_io_imem_req_valid),
    .io_imem_req_bits_addr(fetch_io_imem_req_bits_addr),
    .io_imem_resp_ready(fetch_io_imem_resp_ready),
    .io_imem_resp_valid(fetch_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(fetch_io_imem_resp_bits_rdata)
  );
  ysyx_210340_CacheController icache ( // @[Core.scala 20:22]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_sram0_cen(icache_io_sram0_cen), 
    .io_sram0_wen(icache_io_sram0_wen), 
    .io_sram0_addr(icache_io_sram0_addr), 
    .io_sram0_wdata(icache_io_sram0_wdata), 
    .io_sram0_rdata(icache_io_sram0_rdata), 
    .io_sram1_cen(icache_io_sram1_cen), 
    .io_sram1_wen(icache_io_sram1_wen), 
    .io_sram1_addr(icache_io_sram1_addr), 
    .io_sram1_wdata(icache_io_sram1_wdata), 
    .io_sram1_rdata(icache_io_sram1_rdata),  
    .io_sram2_cen(icache_io_sram2_cen), 
    .io_sram2_wen(icache_io_sram2_wen), 
    .io_sram2_addr(icache_io_sram2_addr), 
    .io_sram2_wdata(icache_io_sram2_wdata), 
    .io_sram2_rdata(icache_io_sram2_rdata),   
    .io_sram3_cen(icache_io_sram3_cen), 
    .io_sram3_wen(icache_io_sram3_wen), 
    .io_sram3_addr(icache_io_sram3_addr), 
    .io_sram3_wdata(icache_io_sram3_wdata), 
    .io_sram3_rdata(icache_io_sram3_rdata),   
    .io_in_req_ready(icache_io_in_req_ready),
    .io_in_req_valid(icache_io_in_req_valid),
    .io_in_req_bits_addr(icache_io_in_req_bits_addr),
    .io_in_resp_ready(icache_io_in_resp_ready),
    .io_in_resp_valid(icache_io_in_resp_valid),
    .io_in_resp_bits_rdata(icache_io_in_resp_bits_rdata),
    .io_out_cache_req_ready(icache_io_out_cache_req_ready),
    .io_out_cache_req_valid(icache_io_out_cache_req_valid),
    .io_out_cache_req_bits_addr(icache_io_out_cache_req_bits_addr),
    .io_out_cache_req_bits_aen(icache_io_out_cache_req_bits_aen),
    .io_out_cache_req_bits_ren(icache_io_out_cache_req_bits_ren),
    .io_out_cache_req_bits_wdata(icache_io_out_cache_req_bits_wdata),
    .io_out_cache_req_bits_wlast(icache_io_out_cache_req_bits_wlast),
    .io_out_cache_req_bits_wen(icache_io_out_cache_req_bits_wen),
    .io_out_cache_resp_ready(icache_io_out_cache_resp_ready),
    .io_out_cache_resp_valid(icache_io_out_cache_resp_valid),
    .io_out_cache_resp_bits_rdata(icache_io_out_cache_resp_bits_rdata),
    .io_out_cache_resp_bits_rlast(icache_io_out_cache_resp_bits_rlast),
    .io_out_uncache_req_ready(icache_io_out_uncache_req_ready),
    .io_out_uncache_req_valid(icache_io_out_uncache_req_valid),
    .io_out_uncache_req_bits_addr(icache_io_out_uncache_req_bits_addr),
    .io_out_uncache_req_bits_ren(icache_io_out_uncache_req_bits_ren),
    .io_out_uncache_req_bits_wdata(icache_io_out_uncache_req_bits_wdata),
    .io_out_uncache_req_bits_wmask(icache_io_out_uncache_req_bits_wmask),
    .io_out_uncache_req_bits_wen(icache_io_out_uncache_req_bits_wen),
    .io_out_uncache_req_bits_size(icache_io_out_uncache_req_bits_size),
    .io_out_uncache_resp_ready(icache_io_out_uncache_resp_ready),
    .io_out_uncache_resp_valid(icache_io_out_uncache_resp_valid),
    .io_out_uncache_resp_bits_rdata(icache_io_out_uncache_resp_bits_rdata),
    .fence_i(icache_fence_i),
    .dcache_fi_complete(icache_dcache_fi_complete)
  );
  ysyx_210340_PipelineReg if_id_reg ( // @[Core.scala 25:25]
    .clock(if_id_reg_clock),
    .reset(if_id_reg_reset),
    .io_in_pc(if_id_reg_io_in_pc),
    .io_in_inst(if_id_reg_io_in_inst),
    .io_in_imem_hs(if_id_reg_io_in_imem_hs),
    .io_out_pc(if_id_reg_io_out_pc),
    .io_out_inst(if_id_reg_io_out_inst),
    .io_out_imem_hs(if_id_reg_io_out_imem_hs),
    .io_flush(if_id_reg_io_flush),
    .io_stall(if_id_reg_io_stall)
  );
  ysyx_210340_Decode decode ( // @[Core.scala 30:22]
    .io_inst(decode_io_inst),
    .io_rs1_addr(decode_io_rs1_addr),
    .io_rs1_type(decode_io_rs1_type),
    .io_rs2_addr(decode_io_rs2_addr),
    .io_rs2_type(decode_io_rs2_type),
    .io_rd_addr(decode_io_rd_addr),
    .io_rd_en(decode_io_rd_en),
    .io_op_type(decode_io_op_type),
    .io_fuType(decode_io_fuType),
    .io_imm(decode_io_imm),
    .io_csr_imm(decode_io_csr_imm)
  );
  ysyx_210340_RegFile rf ( // @[Core.scala 33:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_pc(rf_io_pc),
    .io_rs1_addr(rf_io_rs1_addr),
    .io_rs2_addr(rf_io_rs2_addr),
    .io_rs1_type(rf_io_rs1_type),
    .io_rs2_type(rf_io_rs2_type),
    .io_rd_addr(rf_io_rd_addr),
    .io_rd_en(rf_io_rd_en),
    .io_rd_data(rf_io_rd_data),
    .io_imm(rf_io_imm),
    .io_csr_imm(rf_io_csr_imm),
    .io_irq(rf_io_irq),
    .io_rs1(rf_io_rs1),
    .io_rs2(rf_io_rs2),
    .io_src2(rf_io_src2)
  );
  ysyx_210340_Execution execution ( // @[Core.scala 42:25]
    .io_pc(execution_io_pc),
    .io_op_type(execution_io_op_type),
    .io_rs1(execution_io_rs1),
    .io_rs2(execution_io_rs2),
    .io_src2(execution_io_src2),
    .io_fuType(execution_io_fuType),
    .io_imm(execution_io_imm),
    .io_csr_Jmp_addr(execution_io_csr_Jmp_addr),
    .io_csr_Jmp_en(execution_io_csr_Jmp_en),
    .io_csr_data(execution_io_csr_data),
    .io_br_en(execution_io_br_en),
    .io_br_addr(execution_io_br_addr),
    .io_rd_data(execution_io_rd_data),
    .fence_i_0(execution_fence_i_0)
  );
  ysyx_210340_PipelineReg_1 id_ex_reg ( // @[Core.scala 49:25]
    .clock(id_ex_reg_clock),
    .reset(id_ex_reg_reset),
    .io_in_pc(id_ex_reg_io_in_pc),
    .io_in_br_en(id_ex_reg_io_in_br_en),
    .io_in_br_addr(id_ex_reg_io_in_br_addr),
    .io_in_op_type(id_ex_reg_io_in_op_type),
    .io_in_fuType(id_ex_reg_io_in_fuType),
    .io_in_rs1(id_ex_reg_io_in_rs1),
    .io_in_rs2(id_ex_reg_io_in_rs2),
    .io_in_rd_addr(id_ex_reg_io_in_rd_addr),
    .io_in_src2(id_ex_reg_io_in_src2),
    .io_in_rd_en(id_ex_reg_io_in_rd_en),
    .io_in_imem_hs(id_ex_reg_io_in_imem_hs),
    .io_in_rd_data(id_ex_reg_io_in_rd_data),
    .io_out_pc(id_ex_reg_io_out_pc),
    .io_out_br_en(id_ex_reg_io_out_br_en),
    .io_out_br_addr(id_ex_reg_io_out_br_addr),
    .io_out_op_type(id_ex_reg_io_out_op_type),
    .io_out_fuType(id_ex_reg_io_out_fuType),
    .io_out_rs1(id_ex_reg_io_out_rs1),
    .io_out_rs2(id_ex_reg_io_out_rs2),
    .io_out_rd_addr(id_ex_reg_io_out_rd_addr),
    .io_out_src2(id_ex_reg_io_out_src2),
    .io_out_rd_en(id_ex_reg_io_out_rd_en),
    .io_out_imem_hs(id_ex_reg_io_out_imem_hs),
    .io_out_rd_data(id_ex_reg_io_out_rd_data),
    .io_stall(id_ex_reg_io_stall)
  );
  ysyx_210340_Mem mem ( // @[Core.scala 67:19]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_pc(mem_io_pc),
    .io_op_type(mem_io_op_type),
    .io_rs1(mem_io_rs1),
    .io_rs2(mem_io_rs2),
    .io_src2(mem_io_src2),
    .io_fuType(mem_io_fuType),
    .io_irq(mem_io_irq),
    .io_mem_en(mem_io_mem_en),
    .io_rd_data(mem_io_rd_data),
    .io_busy(mem_io_busy),
    .io_dmem_hs(mem_io_dmem_hs),
    .io_resp_success(mem_io_resp_success),
    .io_dmem_req_ready(mem_io_dmem_req_ready),
    .io_dmem_req_valid(mem_io_dmem_req_valid),
    .io_dmem_req_bits_addr(mem_io_dmem_req_bits_addr),
    .io_dmem_req_bits_ren(mem_io_dmem_req_bits_ren),
    .io_dmem_req_bits_wdata(mem_io_dmem_req_bits_wdata),
    .io_dmem_req_bits_wmask(mem_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wen(mem_io_dmem_req_bits_wen),
    .io_dmem_req_bits_size(mem_io_dmem_req_bits_size),
    .io_dmem_resp_ready(mem_io_dmem_resp_ready),
    .io_dmem_resp_valid(mem_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(mem_io_dmem_resp_bits_rdata)
  );
  ysyx_210340_CSR csr ( // @[Core.scala 77:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_pc(csr_io_pc),
    .io_fuType(csr_io_fuType),
    .io_op_type(csr_io_op_type),
    .io_rs1(csr_io_rs1),
    .io_rs2(csr_io_rs2),
    .io_if_valid(csr_io_if_valid),
    .io_mem_en(csr_io_mem_en),
    .io_mem_valid(csr_io_mem_valid),
    .io_csr_Jmp_addr(csr_io_csr_Jmp_addr),
    .io_csr_Jmp_en(csr_io_csr_Jmp_en),
    .io_csr_data(csr_io_csr_data),
    .io_irq(csr_io_irq),
    .mtip_0(csr_mtip_0)
  );
  ysyx_210340_CacheBusCrossbar1to2 crossbar1to2 ( // @[Core.scala 87:28]
    .clock(crossbar1to2_clock),
    .io_in_req_ready(crossbar1to2_io_in_req_ready),
    .io_in_req_valid(crossbar1to2_io_in_req_valid),
    .io_in_req_bits_addr(crossbar1to2_io_in_req_bits_addr),
    .io_in_req_bits_ren(crossbar1to2_io_in_req_bits_ren),
    .io_in_req_bits_wdata(crossbar1to2_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(crossbar1to2_io_in_req_bits_wmask),
    .io_in_req_bits_wen(crossbar1to2_io_in_req_bits_wen),
    .io_in_req_bits_size(crossbar1to2_io_in_req_bits_size),
    .io_in_resp_ready(crossbar1to2_io_in_resp_ready),
    .io_in_resp_valid(crossbar1to2_io_in_resp_valid),
    .io_in_resp_bits_rdata(crossbar1to2_io_in_resp_bits_rdata),
    .io_out_0_req_ready(crossbar1to2_io_out_0_req_ready),
    .io_out_0_req_valid(crossbar1to2_io_out_0_req_valid),
    .io_out_0_req_bits_addr(crossbar1to2_io_out_0_req_bits_addr),
    .io_out_0_req_bits_ren(crossbar1to2_io_out_0_req_bits_ren),
    .io_out_0_req_bits_wdata(crossbar1to2_io_out_0_req_bits_wdata),
    .io_out_0_req_bits_wmask(crossbar1to2_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wen(crossbar1to2_io_out_0_req_bits_wen),
    .io_out_0_req_bits_size(crossbar1to2_io_out_0_req_bits_size),
    .io_out_0_resp_ready(crossbar1to2_io_out_0_resp_ready),
    .io_out_0_resp_valid(crossbar1to2_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(crossbar1to2_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(crossbar1to2_io_out_1_req_ready),
    .io_out_1_req_valid(crossbar1to2_io_out_1_req_valid),
    .io_out_1_req_bits_addr(crossbar1to2_io_out_1_req_bits_addr),
    .io_out_1_req_bits_ren(crossbar1to2_io_out_1_req_bits_ren),
    .io_out_1_req_bits_wdata(crossbar1to2_io_out_1_req_bits_wdata),
    .io_out_1_req_bits_wmask(crossbar1to2_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wen(crossbar1to2_io_out_1_req_bits_wen),
    .io_out_1_req_bits_size(crossbar1to2_io_out_1_req_bits_size),
    .io_out_1_resp_ready(crossbar1to2_io_out_1_resp_ready),
    .io_out_1_resp_valid(crossbar1to2_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(crossbar1to2_io_out_1_resp_bits_rdata),
    .io_to_1(crossbar1to2_io_to_1)
  );
  ysyx_210340_CacheController_1 dcache ( // @[Core.scala 94:22]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_sram4_cen(dcache_io_sram4_cen), 
    .io_sram4_wen(dcache_io_sram4_wen), 
    .io_sram4_addr(dcache_io_sram4_addr), 
    .io_sram4_wdata(dcache_io_sram4_wdata), 
    .io_sram4_rdata(dcache_io_sram4_rdata), 
    .io_sram5_cen(dcache_io_sram5_cen), 
    .io_sram5_wen(dcache_io_sram5_wen), 
    .io_sram5_addr(dcache_io_sram5_addr), 
    .io_sram5_wdata(dcache_io_sram5_wdata), 
    .io_sram5_rdata(dcache_io_sram5_rdata), 
    .io_sram6_cen(dcache_io_sram6_cen), 
    .io_sram6_wen(dcache_io_sram6_wen), 
    .io_sram6_addr(dcache_io_sram6_addr), 
    .io_sram6_wdata(dcache_io_sram6_wdata), 
    .io_sram6_rdata(dcache_io_sram6_rdata),   
    .io_sram7_cen(dcache_io_sram7_cen), 
    .io_sram7_wen(dcache_io_sram7_wen), 
    .io_sram7_addr(dcache_io_sram7_addr), 
    .io_sram7_wdata(dcache_io_sram7_wdata), 
    .io_sram7_rdata(dcache_io_sram7_rdata),  
    .io_in_req_ready(dcache_io_in_req_ready),
    .io_in_req_valid(dcache_io_in_req_valid),
    .io_in_req_bits_addr(dcache_io_in_req_bits_addr),
    .io_in_req_bits_ren(dcache_io_in_req_bits_ren),
    .io_in_req_bits_wdata(dcache_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(dcache_io_in_req_bits_wmask),
    .io_in_req_bits_wen(dcache_io_in_req_bits_wen),
    .io_in_req_bits_size(dcache_io_in_req_bits_size),
    .io_in_resp_ready(dcache_io_in_resp_ready),
    .io_in_resp_valid(dcache_io_in_resp_valid),
    .io_in_resp_bits_rdata(dcache_io_in_resp_bits_rdata),
    .io_out_cache_req_ready(dcache_io_out_cache_req_ready),
    .io_out_cache_req_valid(dcache_io_out_cache_req_valid),
    .io_out_cache_req_bits_addr(dcache_io_out_cache_req_bits_addr),
    .io_out_cache_req_bits_aen(dcache_io_out_cache_req_bits_aen),
    .io_out_cache_req_bits_ren(dcache_io_out_cache_req_bits_ren),
    .io_out_cache_req_bits_wdata(dcache_io_out_cache_req_bits_wdata),
    .io_out_cache_req_bits_wlast(dcache_io_out_cache_req_bits_wlast),
    .io_out_cache_req_bits_wen(dcache_io_out_cache_req_bits_wen),
    .io_out_cache_resp_ready(dcache_io_out_cache_resp_ready),
    .io_out_cache_resp_valid(dcache_io_out_cache_resp_valid),
    .io_out_cache_resp_bits_rdata(dcache_io_out_cache_resp_bits_rdata),
    .io_out_cache_resp_bits_rlast(dcache_io_out_cache_resp_bits_rlast),
    .io_out_uncache_req_ready(dcache_io_out_uncache_req_ready),
    .io_out_uncache_req_valid(dcache_io_out_uncache_req_valid),
    .io_out_uncache_req_bits_addr(dcache_io_out_uncache_req_bits_addr),
    .io_out_uncache_req_bits_ren(dcache_io_out_uncache_req_bits_ren),
    .io_out_uncache_req_bits_wdata(dcache_io_out_uncache_req_bits_wdata),
    .io_out_uncache_req_bits_wmask(dcache_io_out_uncache_req_bits_wmask),
    .io_out_uncache_req_bits_wen(dcache_io_out_uncache_req_bits_wen),
    .io_out_uncache_req_bits_size(dcache_io_out_uncache_req_bits_size),
    .io_out_uncache_resp_ready(dcache_io_out_uncache_resp_ready),
    .io_out_uncache_resp_valid(dcache_io_out_uncache_resp_valid),
    .io_out_uncache_resp_bits_rdata(dcache_io_out_uncache_resp_bits_rdata),
    .fence_i(dcache_fence_i),
    .dcache_fi_complete(dcache_dcache_fi_complete)
  );

  assign io_sram0_addr = icache_io_sram0_addr; // @[cpu.scala 163:22]
  assign io_sram0_cen = icache_io_sram0_cen; // @[cpu.scala 163:22]
  assign io_sram0_wen = icache_io_sram0_wen; // @[cpu.scala 163:22]
  assign io_sram0_wdata = icache_io_sram0_wdata; // @[cpu.scala 163:22]
  assign io_sram1_addr = icache_io_sram1_addr; // @[cpu.scala 164:22]
  assign io_sram1_cen = icache_io_sram1_cen; // @[cpu.scala 164:22]
  assign io_sram1_wen = icache_io_sram1_wen; // @[cpu.scala 164:22]
  assign io_sram1_wdata = icache_io_sram1_wdata; // @[cpu.scala 164:22]
  assign io_sram2_addr = icache_io_sram2_addr; // @[cpu.scala 165:22]
  assign io_sram2_cen = icache_io_sram2_cen; // @[cpu.scala 165:22]
  assign io_sram2_wen = icache_io_sram2_wen; // @[cpu.scala 165:22]
  assign io_sram2_wdata = icache_io_sram2_wdata; // @[cpu.scala 165:22]
  assign io_sram3_addr = icache_io_sram3_addr; // @[cpu.scala 166:22]
  assign io_sram3_cen = icache_io_sram3_cen; // @[cpu.scala 166:22]
  assign io_sram3_wen = icache_io_sram3_wen; // @[cpu.scala 166:22]
  assign io_sram3_wdata = icache_io_sram3_wdata; // @[cpu.scala 166:22]
  assign io_sram4_addr = dcache_io_sram4_addr; // @[cpu.scala 167:22]
  assign io_sram4_cen = dcache_io_sram4_cen; // @[cpu.scala 167:22]
  assign io_sram4_wen = dcache_io_sram4_wen; // @[cpu.scala 167:22]
  assign io_sram4_wdata = dcache_io_sram4_wdata; // @[cpu.scala 167:22]
  assign io_sram5_addr = dcache_io_sram5_addr; // @[cpu.scala 168:22]
  assign io_sram5_cen = dcache_io_sram5_cen; // @[cpu.scala 168:22]
  assign io_sram5_wen = dcache_io_sram5_wen; // @[cpu.scala 168:22]
  assign io_sram5_wdata = dcache_io_sram5_wdata; // @[cpu.scala 168:22]
  assign io_sram6_addr = dcache_io_sram6_addr; // @[cpu.scala 169:22]
  assign io_sram6_cen = dcache_io_sram6_cen; // @[cpu.scala 169:22]
  assign io_sram6_wen = dcache_io_sram6_wen; // @[cpu.scala 169:22]
  assign io_sram6_wdata = dcache_io_sram6_wdata; // @[cpu.scala 169:22]
  assign io_sram7_addr = dcache_io_sram7_addr; // @[cpu.scala 170:22]
  assign io_sram7_cen = dcache_io_sram7_cen; // @[cpu.scala 170:22]
  assign io_sram7_wen = dcache_io_sram7_wen; // @[cpu.scala 170:22]
  assign io_sram7_wdata = dcache_io_sram7_wdata; // @[cpu.scala 170:22]

  assign icache_io_sram0_rdata = io_sram0_rdata;
  assign icache_io_sram1_rdata = io_sram1_rdata;
  assign icache_io_sram2_rdata = io_sram2_rdata;
  assign icache_io_sram3_rdata = io_sram3_rdata;
  assign dcache_io_sram4_rdata = io_sram4_rdata;
  assign dcache_io_sram5_rdata = io_sram5_rdata;
  assign dcache_io_sram6_rdata = io_sram6_rdata;
  assign dcache_io_sram7_rdata = io_sram7_rdata;


  ysyx_210340_Clint clint ( // @[Core.scala 99:21]
    .clock(clint_clock),
    .reset(clint_reset),
    .io_in_req_ready(clint_io_in_req_ready),
    .io_in_req_valid(clint_io_in_req_valid),
    .io_in_req_bits_addr(clint_io_in_req_bits_addr),
    .io_in_req_bits_ren(clint_io_in_req_bits_ren),
    .io_in_req_bits_wdata(clint_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(clint_io_in_req_bits_wmask),
    .io_in_req_bits_wen(clint_io_in_req_bits_wen),
    .io_in_resp_ready(clint_io_in_resp_ready),
    .io_in_resp_valid(clint_io_in_resp_valid),
    .io_in_resp_bits_rdata(clint_io_in_resp_bits_rdata),
    .mtip_0(clint_mtip_0)
  );
  assign io_core_bus_0_req_valid = icache_io_out_cache_req_valid; // @[Core.scala 22:23]
  assign io_core_bus_0_req_bits_addr = icache_io_out_cache_req_bits_addr; // @[Core.scala 22:23]
  assign io_core_bus_0_req_bits_aen = icache_io_out_cache_req_bits_aen; // @[Core.scala 22:23]
  assign io_core_bus_0_req_bits_ren = icache_io_out_cache_req_bits_ren; // @[Core.scala 22:23]
  assign io_core_bus_0_req_bits_wdata = icache_io_out_cache_req_bits_wdata; // @[Core.scala 22:23]
  assign io_core_bus_0_req_bits_wlast = icache_io_out_cache_req_bits_wlast; // @[Core.scala 22:23]
  assign io_core_bus_0_req_bits_wen = icache_io_out_cache_req_bits_wen; // @[Core.scala 22:23]
  assign io_core_bus_0_resp_ready = icache_io_out_cache_resp_ready; // @[Core.scala 22:23]
  assign io_core_bus_1_req_valid = dcache_io_out_cache_req_valid; // @[Core.scala 96:23]
  assign io_core_bus_1_req_bits_addr = dcache_io_out_cache_req_bits_addr; // @[Core.scala 96:23]
  assign io_core_bus_1_req_bits_aen = dcache_io_out_cache_req_bits_aen; // @[Core.scala 96:23]
  assign io_core_bus_1_req_bits_ren = dcache_io_out_cache_req_bits_ren; // @[Core.scala 96:23]
  assign io_core_bus_1_req_bits_wdata = dcache_io_out_cache_req_bits_wdata; // @[Core.scala 96:23]
  assign io_core_bus_1_req_bits_wlast = dcache_io_out_cache_req_bits_wlast; // @[Core.scala 96:23]
  assign io_core_bus_1_req_bits_wen = dcache_io_out_cache_req_bits_wen; // @[Core.scala 96:23]
  assign io_core_bus_1_resp_ready = dcache_io_out_cache_resp_ready; // @[Core.scala 96:23]
  assign io_core_bus_2_req_valid = icache_io_out_uncache_req_valid; // @[Core.scala 23:25]
  assign io_core_bus_2_req_bits_addr = icache_io_out_uncache_req_bits_addr; // @[Core.scala 23:25]
  assign io_core_bus_2_req_bits_ren = icache_io_out_uncache_req_bits_ren; // @[Core.scala 23:25]
  assign io_core_bus_2_req_bits_wdata = icache_io_out_uncache_req_bits_wdata; // @[Core.scala 23:25]
  assign io_core_bus_2_req_bits_wmask = icache_io_out_uncache_req_bits_wmask; // @[Core.scala 23:25]
  assign io_core_bus_2_req_bits_wen = icache_io_out_uncache_req_bits_wen; // @[Core.scala 23:25]
  assign io_core_bus_2_req_bits_size = icache_io_out_uncache_req_bits_size; // @[Core.scala 23:25]
  assign io_core_bus_2_resp_ready = icache_io_out_uncache_resp_ready; // @[Core.scala 23:25]
  assign io_core_bus_3_req_valid = dcache_io_out_uncache_req_valid; // @[Core.scala 97:25]
  assign io_core_bus_3_req_bits_addr = dcache_io_out_uncache_req_bits_addr; // @[Core.scala 97:25]
  assign io_core_bus_3_req_bits_ren = dcache_io_out_uncache_req_bits_ren; // @[Core.scala 97:25]
  assign io_core_bus_3_req_bits_wdata = dcache_io_out_uncache_req_bits_wdata; // @[Core.scala 97:25]
  assign io_core_bus_3_req_bits_wmask = dcache_io_out_uncache_req_bits_wmask; // @[Core.scala 97:25]
  assign io_core_bus_3_req_bits_wen = dcache_io_out_uncache_req_bits_wen; // @[Core.scala 97:25]
  assign io_core_bus_3_req_bits_size = dcache_io_out_uncache_req_bits_size; // @[Core.scala 97:25]
  assign io_core_bus_3_resp_ready = dcache_io_out_uncache_resp_ready; // @[Core.scala 97:25]
  assign fetch_clock = clock;
  assign fetch_reset = reset;
  assign fetch_io_stall = mem_io_busy; // @[Core.scala 122:18]
  assign fetch_io_flush = execution_io_br_en | execution_io_csr_Jmp_en; // @[Core.scala 123:40]
  assign fetch_io_br_en = id_ex_reg_io_out_br_en; // @[Core.scala 62:20]
  assign fetch_io_br_addr = id_ex_reg_io_out_br_addr; // @[Core.scala 63:20]
  assign fetch_io_imem_req_ready = icache_io_in_req_ready; // @[Core.scala 21:16]
  assign fetch_io_imem_resp_valid = icache_io_in_resp_valid; // @[Core.scala 21:16]
  assign fetch_io_imem_resp_bits_rdata = icache_io_in_resp_bits_rdata; // @[Core.scala 21:16]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_in_req_valid = fetch_io_imem_req_valid; // @[Core.scala 21:16]
  assign icache_io_in_req_bits_addr = fetch_io_imem_req_bits_addr; // @[Core.scala 21:16]
  assign icache_io_in_resp_ready = fetch_io_imem_resp_ready; // @[Core.scala 21:16]
  assign icache_io_out_cache_req_ready = io_core_bus_0_req_ready; // @[Core.scala 22:23]
  assign icache_io_out_cache_resp_valid = io_core_bus_0_resp_valid; // @[Core.scala 22:23]
  assign icache_io_out_cache_resp_bits_rdata = io_core_bus_0_resp_bits_rdata; // @[Core.scala 22:23]
  assign icache_io_out_cache_resp_bits_rlast = io_core_bus_0_resp_bits_rlast; // @[Core.scala 22:23]
  assign icache_io_out_uncache_req_ready = io_core_bus_2_req_ready; // @[Core.scala 23:25]
  assign icache_io_out_uncache_resp_valid = io_core_bus_2_resp_valid; // @[Core.scala 23:25]
  assign icache_io_out_uncache_resp_bits_rdata = io_core_bus_2_resp_bits_rdata; // @[Core.scala 23:25]
  assign icache_fence_i = execution_fence_i_0;
  assign icache_dcache_fi_complete = dcache_dcache_fi_complete;
  assign if_id_reg_clock = clock;
  assign if_id_reg_reset = reset;
  assign if_id_reg_io_in_pc = fetch_io_out_pc; // @[Core.scala 26:19]
  assign if_id_reg_io_in_inst = fetch_io_out_inst; // @[Core.scala 26:19]
  assign if_id_reg_io_in_imem_hs = fetch_io_out_imem_hs; // @[Core.scala 26:19]
  assign if_id_reg_io_flush = execution_io_br_en | execution_io_csr_Jmp_en; // @[Core.scala 127:45]
  assign if_id_reg_io_stall = mem_io_busy; // @[Core.scala 126:23]
  assign decode_io_inst = if_id_reg_io_out_inst; // @[Core.scala 31:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_pc = if_id_reg_io_out_pc; // @[Core.scala 34:18]
  assign rf_io_rs1_addr = decode_io_rs1_addr; // @[Core.scala 35:18]
  assign rf_io_rs2_addr = decode_io_rs2_addr; // @[Core.scala 36:18]
  assign rf_io_rs1_type = decode_io_rs1_type; // @[Core.scala 37:18]
  assign rf_io_rs2_type = decode_io_rs2_type; // @[Core.scala 38:18]
  assign rf_io_rd_addr = id_ex_reg_io_out_rd_addr; // @[Core.scala 109:29]
  assign rf_io_rd_en = mem_io_mem_en & ~id_ex_reg_io_out_op_type[3] ? reg_wen_REG : id_ex_reg_io_out_rd_en; // @[Core.scala 75:20]
  assign rf_io_rd_data = csr_io_fuType == 3'h3 ? execution_io_csr_data : _rf_io_rd_data_T_4; // @[Core.scala 108:35]
  assign rf_io_imm = decode_io_imm; // @[Core.scala 39:18]
  assign rf_io_csr_imm = decode_io_csr_imm; // @[Core.scala 40:18]
  assign rf_io_irq = csr_io_irq; // @[Core.scala 106:29]
  assign execution_io_pc = if_id_reg_io_out_pc; // @[Core.scala 43:24]
  assign execution_io_op_type = decode_io_op_type; // @[Core.scala 44:24]
  assign execution_io_rs1 = rf_io_rs1; // @[Core.scala 112:24]
  assign execution_io_rs2 = rf_io_rs2; // @[Core.scala 113:24]
  assign execution_io_src2 = rf_io_src2; // @[Core.scala 114:24]
  assign execution_io_fuType = decode_io_fuType; // @[Core.scala 45:24]
  assign execution_io_imm = decode_io_imm; // @[Core.scala 47:24]
  assign execution_io_csr_Jmp_addr = csr_io_csr_Jmp_addr; // @[Core.scala 102:29]
  assign execution_io_csr_Jmp_en = csr_io_csr_Jmp_en; // @[Core.scala 103:29]
  assign execution_io_csr_data = csr_io_csr_data; // @[Core.scala 104:29]
  assign id_ex_reg_clock = clock;
  assign id_ex_reg_reset = reset;
  assign id_ex_reg_io_in_pc = if_id_reg_io_out_pc; // @[Core.scala 54:27]
  assign id_ex_reg_io_in_br_en = execution_io_br_en; // @[Core.scala 50:27]
  assign id_ex_reg_io_in_br_addr = execution_io_br_addr; // @[Core.scala 51:27]
  assign id_ex_reg_io_in_op_type = decode_io_op_type; // @[Core.scala 52:27]
  assign id_ex_reg_io_in_fuType = decode_io_fuType; // @[Core.scala 53:27]
  assign id_ex_reg_io_in_rs1 = rf_io_rs1; // @[Core.scala 116:24]
  assign id_ex_reg_io_in_rs2 = rf_io_rs2; // @[Core.scala 117:24]
  assign id_ex_reg_io_in_rd_addr = decode_io_rd_addr; // @[Core.scala 56:27]
  assign id_ex_reg_io_in_src2 = rf_io_src2; // @[Core.scala 115:24]
  assign id_ex_reg_io_in_rd_en = decode_io_rd_en; // @[Core.scala 58:27]
  assign id_ex_reg_io_in_imem_hs = if_id_reg_io_out_imem_hs; // @[Core.scala 59:27]
  assign id_ex_reg_io_in_rd_data = execution_io_rd_data; // @[Core.scala 60:27]
  assign id_ex_reg_io_stall = mem_io_busy; // @[Core.scala 129:23]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_pc = id_ex_reg_io_out_pc; // @[Core.scala 68:18]
  assign mem_io_op_type = id_ex_reg_io_out_op_type; // @[Core.scala 69:18]
  assign mem_io_rs1 = id_ex_reg_io_out_rs1; // @[Core.scala 71:18]
  assign mem_io_rs2 = id_ex_reg_io_out_rs2; // @[Core.scala 72:18]
  assign mem_io_src2 = id_ex_reg_io_out_src2; // @[Core.scala 73:18]
  assign mem_io_fuType = id_ex_reg_io_out_fuType; // @[Core.scala 70:18]
  assign mem_io_irq = csr_io_irq; // @[Core.scala 110:29]
  assign mem_io_dmem_req_ready = crossbar1to2_io_in_req_ready; // @[Core.scala 88:22]
  assign mem_io_dmem_resp_valid = crossbar1to2_io_in_resp_valid; // @[Core.scala 88:22]
  assign mem_io_dmem_resp_bits_rdata = crossbar1to2_io_in_resp_bits_rdata; // @[Core.scala 88:22]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_pc = id_ex_reg_io_out_pc; // @[Core.scala 78:20]
  assign csr_io_fuType = id_ex_reg_io_out_fuType; // @[Core.scala 79:20]
  assign csr_io_op_type = id_ex_reg_io_out_op_type; // @[Core.scala 80:20]
  assign csr_io_rs1 = id_ex_reg_io_out_rs1; // @[Core.scala 81:20]
  assign csr_io_rs2 = id_ex_reg_io_out_rs2; // @[Core.scala 82:20]
  assign csr_io_if_valid = id_ex_reg_io_out_imem_hs; // @[Core.scala 83:20]
  assign csr_io_mem_en = mem_io_mem_en; // @[Core.scala 84:20]
  assign csr_io_mem_valid = mem_io_dmem_hs; // @[Core.scala 85:20]
  assign csr_mtip_0 = clint_mtip_0;
  assign crossbar1to2_clock = clock;
  assign crossbar1to2_io_in_req_valid = mem_io_dmem_req_valid; // @[Core.scala 88:22]
  assign crossbar1to2_io_in_req_bits_addr = mem_io_dmem_req_bits_addr; // @[Core.scala 88:22]
  assign crossbar1to2_io_in_req_bits_ren = mem_io_dmem_req_bits_ren; // @[Core.scala 88:22]
  assign crossbar1to2_io_in_req_bits_wdata = mem_io_dmem_req_bits_wdata; // @[Core.scala 88:22]
  assign crossbar1to2_io_in_req_bits_wmask = mem_io_dmem_req_bits_wmask; // @[Core.scala 88:22]
  assign crossbar1to2_io_in_req_bits_wen = mem_io_dmem_req_bits_wen; // @[Core.scala 88:22]
  assign crossbar1to2_io_in_req_bits_size = mem_io_dmem_req_bits_size; // @[Core.scala 88:22]
  assign crossbar1to2_io_in_resp_ready = mem_io_dmem_resp_ready; // @[Core.scala 88:22]
  assign crossbar1to2_io_out_0_req_ready = dcache_io_in_req_ready; // @[Core.scala 95:16]
  assign crossbar1to2_io_out_0_resp_valid = dcache_io_in_resp_valid; // @[Core.scala 95:16]
  assign crossbar1to2_io_out_0_resp_bits_rdata = dcache_io_in_resp_bits_rdata; // @[Core.scala 95:16]
  assign crossbar1to2_io_out_1_req_ready = clint_io_in_req_ready; // @[Core.scala 100:15]
  assign crossbar1to2_io_out_1_resp_valid = clint_io_in_resp_valid; // @[Core.scala 100:15]
  assign crossbar1to2_io_out_1_resp_bits_rdata = clint_io_in_resp_bits_rdata; // @[Core.scala 100:15]
  assign crossbar1to2_io_to_1 = crossbar1to2_io_in_req_bits_addr >= 32'h2000000 & crossbar1to2_io_in_req_bits_addr < 32'h2010000
    ; // @[Core.scala 91:55]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_in_req_valid = crossbar1to2_io_out_0_req_valid; // @[Core.scala 95:16]
  assign dcache_io_in_req_bits_addr = crossbar1to2_io_out_0_req_bits_addr; // @[Core.scala 95:16]
  assign dcache_io_in_req_bits_ren = crossbar1to2_io_out_0_req_bits_ren; // @[Core.scala 95:16]
  assign dcache_io_in_req_bits_wdata = crossbar1to2_io_out_0_req_bits_wdata; // @[Core.scala 95:16]
  assign dcache_io_in_req_bits_wmask = crossbar1to2_io_out_0_req_bits_wmask; // @[Core.scala 95:16]
  assign dcache_io_in_req_bits_wen = crossbar1to2_io_out_0_req_bits_wen; // @[Core.scala 95:16]
  assign dcache_io_in_req_bits_size = crossbar1to2_io_out_0_req_bits_size; // @[Core.scala 95:16]
  assign dcache_io_in_resp_ready = crossbar1to2_io_out_0_resp_ready; // @[Core.scala 95:16]
  assign dcache_io_out_cache_req_ready = io_core_bus_1_req_ready; // @[Core.scala 96:23]
  assign dcache_io_out_cache_resp_valid = io_core_bus_1_resp_valid; // @[Core.scala 96:23]
  assign dcache_io_out_cache_resp_bits_rdata = io_core_bus_1_resp_bits_rdata; // @[Core.scala 96:23]
  assign dcache_io_out_cache_resp_bits_rlast = io_core_bus_1_resp_bits_rlast; // @[Core.scala 96:23]
  assign dcache_io_out_uncache_req_ready = io_core_bus_3_req_ready; // @[Core.scala 97:25]
  assign dcache_io_out_uncache_resp_valid = io_core_bus_3_resp_valid; // @[Core.scala 97:25]
  assign dcache_io_out_uncache_resp_bits_rdata = io_core_bus_3_resp_bits_rdata; // @[Core.scala 97:25]
  assign dcache_fence_i = execution_fence_i_0;
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io_in_req_valid = crossbar1to2_io_out_1_req_valid; // @[Core.scala 100:15]
  assign clint_io_in_req_bits_addr = crossbar1to2_io_out_1_req_bits_addr; // @[Core.scala 100:15]
  assign clint_io_in_req_bits_ren = crossbar1to2_io_out_1_req_bits_ren; // @[Core.scala 100:15]
  assign clint_io_in_req_bits_wdata = crossbar1to2_io_out_1_req_bits_wdata; // @[Core.scala 100:15]
  assign clint_io_in_req_bits_wmask = crossbar1to2_io_out_1_req_bits_wmask; // @[Core.scala 100:15]
  assign clint_io_in_req_bits_wen = crossbar1to2_io_out_1_req_bits_wen; // @[Core.scala 100:15]
  assign clint_io_in_resp_ready = crossbar1to2_io_out_1_resp_ready; // @[Core.scala 100:15]
  always @(posedge clock) begin
    reg_wen_REG <= mem_io_resp_success; // @[Core.scala 75:85]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_wen_REG = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210340_RRArbiter_3(
  input         clock,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input         io_in_0_bits_aen,
  input         io_in_0_bits_ren,
  input  [63:0] io_in_0_bits_wdata,
  input         io_in_0_bits_wlast,
  input         io_in_0_bits_wen,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input         io_in_1_bits_aen,
  input         io_in_1_bits_ren,
  input  [63:0] io_in_1_bits_wdata,
  input         io_in_1_bits_wlast,
  input         io_in_1_bits_wen,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_addr,
  input         io_in_2_bits_ren,
  input  [63:0] io_in_2_bits_wdata,
  input  [7:0]  io_in_2_bits_wmask,
  input         io_in_2_bits_wen,
  input  [1:0]  io_in_2_bits_size,
  input         io_in_3_valid,
  input  [31:0] io_in_3_bits_addr,
  input         io_in_3_bits_ren,
  input  [63:0] io_in_3_bits_wdata,
  input  [7:0]  io_in_3_bits_wmask,
  input         io_in_3_bits_wen,
  input  [1:0]  io_in_3_bits_size,
  input         io_out_ready,
  output        io_out_valid,
  output [3:0]  io_out_bits_id,
  output [31:0] io_out_bits_addr,
  output        io_out_bits_aen,
  output        io_out_bits_ren,
  output [63:0] io_out_bits_wdata,
  output [7:0]  io_out_bits_wmask,
  output        io_out_bits_wlast,
  output        io_out_bits_wen,
  output [7:0]  io_out_bits_len,
  output [1:0]  io_out_bits_size,
  output [1:0]  io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _GEN_1 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16 Arbiter.scala 41:16]
  wire  _GEN_2 = 2'h2 == io_chosen ? io_in_2_valid : _GEN_1; // @[Arbiter.scala 41:16 Arbiter.scala 41:16]
  wire [1:0] _GEN_6 = 2'h2 == io_chosen ? io_in_2_bits_size : 2'h3; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire [7:0] _GEN_10 = 2'h2 == io_chosen ? 8'h0 : 8'h1; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire  _GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_wen : io_in_0_bits_wen; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire  _GEN_14 = 2'h2 == io_chosen ? io_in_2_bits_wen : _GEN_13; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire  _GEN_17 = 2'h1 == io_chosen ? io_in_1_bits_wlast : io_in_0_bits_wlast; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire [7:0] _GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_wmask : 8'hff; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire [63:0] _GEN_25 = 2'h1 == io_chosen ? io_in_1_bits_wdata : io_in_0_bits_wdata; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire [63:0] _GEN_26 = 2'h2 == io_chosen ? io_in_2_bits_wdata : _GEN_25; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire  _GEN_29 = 2'h1 == io_chosen ? io_in_1_bits_ren : io_in_0_bits_ren; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire  _GEN_30 = 2'h2 == io_chosen ? io_in_2_bits_ren : _GEN_29; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire  _GEN_33 = 2'h1 == io_chosen ? io_in_1_bits_aen : io_in_0_bits_aen; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire [31:0] _GEN_37 = 2'h1 == io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire [31:0] _GEN_38 = 2'h2 == io_chosen ? io_in_2_bits_addr : _GEN_37; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire [3:0] _GEN_41 = 2'h1 == io_chosen ? 4'h2 : 4'h1; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire [3:0] _GEN_42 = 2'h2 == io_chosen ? 4'h3 : _GEN_41; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire  _ctrl_validMask_grantMask_lastGrant_T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg [1:0] lastGrant; // @[Reg.scala 15:16]
  wire  grantMask_1 = 2'h1 > lastGrant; // @[Arbiter.scala 67:49]
  wire  grantMask_2 = 2'h2 > lastGrant; // @[Arbiter.scala 67:49]
  wire  grantMask_3 = 2'h3 > lastGrant; // @[Arbiter.scala 67:49]
  wire  validMask_1 = io_in_1_valid & grantMask_1; // @[Arbiter.scala 68:75]
  wire  validMask_2 = io_in_2_valid & grantMask_2; // @[Arbiter.scala 68:75]
  wire  validMask_3 = io_in_3_valid & grantMask_3; // @[Arbiter.scala 68:75]
  wire [1:0] _GEN_45 = io_in_2_valid ? 2'h2 : 2'h3; // @[Arbiter.scala 77:27 Arbiter.scala 77:36]
  wire [1:0] _GEN_46 = io_in_1_valid ? 2'h1 : _GEN_45; // @[Arbiter.scala 77:27 Arbiter.scala 77:36]
  wire [1:0] _GEN_47 = io_in_0_valid ? 2'h0 : _GEN_46; // @[Arbiter.scala 77:27 Arbiter.scala 77:36]
  wire [1:0] _GEN_48 = validMask_3 ? 2'h3 : _GEN_47; // @[Arbiter.scala 79:25 Arbiter.scala 79:34]
  wire [1:0] _GEN_49 = validMask_2 ? 2'h2 : _GEN_48; // @[Arbiter.scala 79:25 Arbiter.scala 79:34]
  assign io_out_valid = 2'h3 == io_chosen ? io_in_3_valid : _GEN_2; // @[Arbiter.scala 41:16 Arbiter.scala 41:16]
  assign io_out_bits_id = 2'h3 == io_chosen ? 4'h4 : _GEN_42; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_out_bits_addr = 2'h3 == io_chosen ? io_in_3_bits_addr : _GEN_38; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_out_bits_aen = 2'h3 == io_chosen | (2'h2 == io_chosen | _GEN_33); // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_out_bits_ren = 2'h3 == io_chosen ? io_in_3_bits_ren : _GEN_30; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_out_bits_wdata = 2'h3 == io_chosen ? io_in_3_bits_wdata : _GEN_26; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_out_bits_wmask = 2'h3 == io_chosen ? io_in_3_bits_wmask : _GEN_22; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_out_bits_wlast = 2'h3 == io_chosen | (2'h2 == io_chosen | _GEN_17); // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_out_bits_wen = 2'h3 == io_chosen ? io_in_3_bits_wen : _GEN_14; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_out_bits_len = 2'h3 == io_chosen ? 8'h0 : _GEN_10; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_out_bits_size = 2'h3 == io_chosen ? io_in_3_bits_size : _GEN_6; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_chosen = validMask_1 ? 2'h1 : _GEN_49; // @[Arbiter.scala 79:25 Arbiter.scala 79:34]
  always @(posedge clock) begin
    if (_ctrl_validMask_grantMask_lastGrant_T) begin // @[Reg.scala 16:19]
      lastGrant <= io_chosen; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lastGrant = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210340_CoreBusCrossbarNto1(
  input         clock,
  output        io_in_0_req_ready,
  input         io_in_0_req_valid,
  input  [31:0] io_in_0_req_bits_addr,
  input         io_in_0_req_bits_aen,
  input         io_in_0_req_bits_ren,
  input  [63:0] io_in_0_req_bits_wdata,
  input         io_in_0_req_bits_wlast,
  input         io_in_0_req_bits_wen,
  input         io_in_0_resp_ready,
  output        io_in_0_resp_valid,
  output [63:0] io_in_0_resp_bits_rdata,
  output        io_in_0_resp_bits_rlast,
  output        io_in_1_req_ready,
  input         io_in_1_req_valid,
  input  [31:0] io_in_1_req_bits_addr,
  input         io_in_1_req_bits_aen,
  input         io_in_1_req_bits_ren,
  input  [63:0] io_in_1_req_bits_wdata,
  input         io_in_1_req_bits_wlast,
  input         io_in_1_req_bits_wen,
  input         io_in_1_resp_ready,
  output        io_in_1_resp_valid,
  output [63:0] io_in_1_resp_bits_rdata,
  output        io_in_1_resp_bits_rlast,
  output        io_in_2_req_ready,
  input         io_in_2_req_valid,
  input  [31:0] io_in_2_req_bits_addr,
  input         io_in_2_req_bits_ren,
  input  [63:0] io_in_2_req_bits_wdata,
  input  [7:0]  io_in_2_req_bits_wmask,
  input         io_in_2_req_bits_wen,
  input  [1:0]  io_in_2_req_bits_size,
  input         io_in_2_resp_ready,
  output        io_in_2_resp_valid,
  output [63:0] io_in_2_resp_bits_rdata,
  output        io_in_3_req_ready,
  input         io_in_3_req_valid,
  input  [31:0] io_in_3_req_bits_addr,
  input         io_in_3_req_bits_ren,
  input  [63:0] io_in_3_req_bits_wdata,
  input  [7:0]  io_in_3_req_bits_wmask,
  input         io_in_3_req_bits_wen,
  input  [1:0]  io_in_3_req_bits_size,
  input         io_in_3_resp_ready,
  output        io_in_3_resp_valid,
  output [63:0] io_in_3_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [3:0]  io_out_req_bits_id,
  output [31:0] io_out_req_bits_addr,
  output        io_out_req_bits_aen,
  output        io_out_req_bits_ren,
  output [63:0] io_out_req_bits_wdata,
  output [7:0]  io_out_req_bits_wmask,
  output        io_out_req_bits_wlast,
  output        io_out_req_bits_wen,
  output [7:0]  io_out_req_bits_len,
  output [1:0]  io_out_req_bits_size,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_id,
  input  [63:0] io_out_resp_bits_rdata,
  input         io_out_resp_bits_rlast
);
  wire  arbiter_clock; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_0_valid; // @[Crossbar.scala 12:23]
  wire [31:0] arbiter_io_in_0_bits_addr; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_0_bits_aen; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_0_bits_ren; // @[Crossbar.scala 12:23]
  wire [63:0] arbiter_io_in_0_bits_wdata; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_0_bits_wlast; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_0_bits_wen; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_1_valid; // @[Crossbar.scala 12:23]
  wire [31:0] arbiter_io_in_1_bits_addr; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_1_bits_aen; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_1_bits_ren; // @[Crossbar.scala 12:23]
  wire [63:0] arbiter_io_in_1_bits_wdata; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_1_bits_wlast; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_1_bits_wen; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_2_valid; // @[Crossbar.scala 12:23]
  wire [31:0] arbiter_io_in_2_bits_addr; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_2_bits_ren; // @[Crossbar.scala 12:23]
  wire [63:0] arbiter_io_in_2_bits_wdata; // @[Crossbar.scala 12:23]
  wire [7:0] arbiter_io_in_2_bits_wmask; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_2_bits_wen; // @[Crossbar.scala 12:23]
  wire [1:0] arbiter_io_in_2_bits_size; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_3_valid; // @[Crossbar.scala 12:23]
  wire [31:0] arbiter_io_in_3_bits_addr; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_3_bits_ren; // @[Crossbar.scala 12:23]
  wire [63:0] arbiter_io_in_3_bits_wdata; // @[Crossbar.scala 12:23]
  wire [7:0] arbiter_io_in_3_bits_wmask; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_3_bits_wen; // @[Crossbar.scala 12:23]
  wire [1:0] arbiter_io_in_3_bits_size; // @[Crossbar.scala 12:23]
  wire  arbiter_io_out_ready; // @[Crossbar.scala 12:23]
  wire  arbiter_io_out_valid; // @[Crossbar.scala 12:23]
  wire [3:0] arbiter_io_out_bits_id; // @[Crossbar.scala 12:23]
  wire [31:0] arbiter_io_out_bits_addr; // @[Crossbar.scala 12:23]
  wire  arbiter_io_out_bits_aen; // @[Crossbar.scala 12:23]
  wire  arbiter_io_out_bits_ren; // @[Crossbar.scala 12:23]
  wire [63:0] arbiter_io_out_bits_wdata; // @[Crossbar.scala 12:23]
  wire [7:0] arbiter_io_out_bits_wmask; // @[Crossbar.scala 12:23]
  wire  arbiter_io_out_bits_wlast; // @[Crossbar.scala 12:23]
  wire  arbiter_io_out_bits_wen; // @[Crossbar.scala 12:23]
  wire [7:0] arbiter_io_out_bits_len; // @[Crossbar.scala 12:23]
  wire [1:0] arbiter_io_out_bits_size; // @[Crossbar.scala 12:23]
  wire [1:0] arbiter_io_chosen; // @[Crossbar.scala 12:23]
  wire  _GEN_0 = io_out_resp_bits_id == 4'h1 & io_in_0_resp_ready; // @[Crossbar.scala 35:46 Crossbar.scala 36:25 Crossbar.scala 32:23]
  wire  _GEN_2 = io_out_resp_bits_id == 4'h2 ? io_in_1_resp_ready : _GEN_0; // @[Crossbar.scala 35:46 Crossbar.scala 36:25]
  wire  _GEN_4 = io_out_resp_bits_id == 4'h3 ? io_in_2_resp_ready : _GEN_2; // @[Crossbar.scala 35:46 Crossbar.scala 36:25]
  ysyx_210340_RRArbiter_3 arbiter ( // @[Crossbar.scala 12:23]
    .clock(arbiter_clock),
    .io_in_0_valid(arbiter_io_in_0_valid),
    .io_in_0_bits_addr(arbiter_io_in_0_bits_addr),
    .io_in_0_bits_aen(arbiter_io_in_0_bits_aen),
    .io_in_0_bits_ren(arbiter_io_in_0_bits_ren),
    .io_in_0_bits_wdata(arbiter_io_in_0_bits_wdata),
    .io_in_0_bits_wlast(arbiter_io_in_0_bits_wlast),
    .io_in_0_bits_wen(arbiter_io_in_0_bits_wen),
    .io_in_1_valid(arbiter_io_in_1_valid),
    .io_in_1_bits_addr(arbiter_io_in_1_bits_addr),
    .io_in_1_bits_aen(arbiter_io_in_1_bits_aen),
    .io_in_1_bits_ren(arbiter_io_in_1_bits_ren),
    .io_in_1_bits_wdata(arbiter_io_in_1_bits_wdata),
    .io_in_1_bits_wlast(arbiter_io_in_1_bits_wlast),
    .io_in_1_bits_wen(arbiter_io_in_1_bits_wen),
    .io_in_2_valid(arbiter_io_in_2_valid),
    .io_in_2_bits_addr(arbiter_io_in_2_bits_addr),
    .io_in_2_bits_ren(arbiter_io_in_2_bits_ren),
    .io_in_2_bits_wdata(arbiter_io_in_2_bits_wdata),
    .io_in_2_bits_wmask(arbiter_io_in_2_bits_wmask),
    .io_in_2_bits_wen(arbiter_io_in_2_bits_wen),
    .io_in_2_bits_size(arbiter_io_in_2_bits_size),
    .io_in_3_valid(arbiter_io_in_3_valid),
    .io_in_3_bits_addr(arbiter_io_in_3_bits_addr),
    .io_in_3_bits_ren(arbiter_io_in_3_bits_ren),
    .io_in_3_bits_wdata(arbiter_io_in_3_bits_wdata),
    .io_in_3_bits_wmask(arbiter_io_in_3_bits_wmask),
    .io_in_3_bits_wen(arbiter_io_in_3_bits_wen),
    .io_in_3_bits_size(arbiter_io_in_3_bits_size),
    .io_out_ready(arbiter_io_out_ready),
    .io_out_valid(arbiter_io_out_valid),
    .io_out_bits_id(arbiter_io_out_bits_id),
    .io_out_bits_addr(arbiter_io_out_bits_addr),
    .io_out_bits_aen(arbiter_io_out_bits_aen),
    .io_out_bits_ren(arbiter_io_out_bits_ren),
    .io_out_bits_wdata(arbiter_io_out_bits_wdata),
    .io_out_bits_wmask(arbiter_io_out_bits_wmask),
    .io_out_bits_wlast(arbiter_io_out_bits_wlast),
    .io_out_bits_wen(arbiter_io_out_bits_wen),
    .io_out_bits_len(arbiter_io_out_bits_len),
    .io_out_bits_size(arbiter_io_out_bits_size),
    .io_chosen(arbiter_io_chosen)
  );
  assign io_in_0_req_ready = arbiter_io_chosen == 2'h0 & io_out_req_ready; // @[Crossbar.scala 20:55]
  assign io_in_0_resp_valid = io_out_resp_bits_id == 4'h1 & io_out_resp_valid; // @[Crossbar.scala 35:46 Crossbar.scala 37:27 Crossbar.scala 31:25]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 30:24]
  assign io_in_0_resp_bits_rlast = io_out_resp_bits_rlast; // @[Crossbar.scala 30:24]
  assign io_in_1_req_ready = arbiter_io_chosen == 2'h1 & io_out_req_ready; // @[Crossbar.scala 20:55]
  assign io_in_1_resp_valid = io_out_resp_bits_id == 4'h2 & io_out_resp_valid; // @[Crossbar.scala 35:46 Crossbar.scala 37:27 Crossbar.scala 31:25]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 30:24]
  assign io_in_1_resp_bits_rlast = io_out_resp_bits_rlast; // @[Crossbar.scala 30:24]
  assign io_in_2_req_ready = arbiter_io_chosen == 2'h2 & io_out_req_ready; // @[Crossbar.scala 20:55]
  assign io_in_2_resp_valid = io_out_resp_bits_id == 4'h3 & io_out_resp_valid; // @[Crossbar.scala 35:46 Crossbar.scala 37:27 Crossbar.scala 31:25]
  assign io_in_2_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 30:24]
  assign io_in_3_req_ready = arbiter_io_chosen == 2'h3 & io_out_req_ready; // @[Crossbar.scala 20:55]
  assign io_in_3_resp_valid = io_out_resp_bits_id == 4'h4 & io_out_resp_valid; // @[Crossbar.scala 35:46 Crossbar.scala 37:27 Crossbar.scala 31:25]
  assign io_in_3_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 30:24]
  assign io_out_req_valid = arbiter_io_out_valid; // @[Crossbar.scala 24:13]
  assign io_out_req_bits_id = arbiter_io_out_bits_id; // @[Crossbar.scala 23:12]
  assign io_out_req_bits_addr = arbiter_io_out_bits_addr; // @[Crossbar.scala 23:12]
  assign io_out_req_bits_aen = arbiter_io_out_bits_aen; // @[Crossbar.scala 23:12]
  assign io_out_req_bits_ren = arbiter_io_out_bits_ren; // @[Crossbar.scala 23:12]
  assign io_out_req_bits_wdata = arbiter_io_out_bits_wdata; // @[Crossbar.scala 23:12]
  assign io_out_req_bits_wmask = arbiter_io_out_bits_wmask; // @[Crossbar.scala 23:12]
  assign io_out_req_bits_wlast = arbiter_io_out_bits_wlast; // @[Crossbar.scala 23:12]
  assign io_out_req_bits_wen = arbiter_io_out_bits_wen; // @[Crossbar.scala 23:12]
  assign io_out_req_bits_len = arbiter_io_out_bits_len; // @[Crossbar.scala 23:12]
  assign io_out_req_bits_size = arbiter_io_out_bits_size; // @[Crossbar.scala 23:12]
  assign io_out_resp_ready = io_out_resp_bits_id == 4'h4 ? io_in_3_resp_ready : _GEN_4; // @[Crossbar.scala 35:46 Crossbar.scala 36:25]
  assign arbiter_clock = clock;
  assign arbiter_io_in_0_valid = io_in_0_req_valid; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_0_bits_aen = io_in_0_req_bits_aen; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_0_bits_ren = io_in_0_req_bits_ren; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_0_bits_wlast = io_in_0_req_bits_wlast; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_0_bits_wen = io_in_0_req_bits_wen; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_1_valid = io_in_1_req_valid; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_1_bits_aen = io_in_1_req_bits_aen; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_1_bits_ren = io_in_1_req_bits_ren; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_1_bits_wlast = io_in_1_req_bits_wlast; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_1_bits_wen = io_in_1_req_bits_wen; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_2_valid = io_in_2_req_valid; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_2_bits_addr = io_in_2_req_bits_addr; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_2_bits_ren = io_in_2_req_bits_ren; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_2_bits_wdata = io_in_2_req_bits_wdata; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_2_bits_wmask = io_in_2_req_bits_wmask; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_2_bits_wen = io_in_2_req_bits_wen; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_2_bits_size = io_in_2_req_bits_size; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_3_valid = io_in_3_req_valid; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_3_bits_addr = io_in_3_req_bits_addr; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_3_bits_ren = io_in_3_req_bits_ren; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_3_bits_wdata = io_in_3_req_bits_wdata; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_3_bits_wmask = io_in_3_req_bits_wmask; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_3_bits_wen = io_in_3_req_bits_wen; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_3_bits_size = io_in_3_req_bits_size; // @[Crossbar.scala 15:22]
  assign arbiter_io_out_ready = io_out_req_ready; // @[Crossbar.scala 25:13]
endmodule
module ysyx_210340_SimpleAxi2Axi(
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [3:0]  io_in_req_bits_id,
  input  [31:0] io_in_req_bits_addr,
  input         io_in_req_bits_aen,
  input         io_in_req_bits_ren,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wlast,
  input         io_in_req_bits_wen,
  input  [7:0]  io_in_req_bits_len,
  input  [1:0]  io_in_req_bits_size,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_id,
  output [63:0] io_in_resp_bits_rdata,
  output        io_in_resp_bits_rlast,
  input         io_out_aw_ready,
  output        io_out_aw_valid,
  output [31:0] io_out_aw_bits_addr,
  output [3:0]  io_out_aw_bits_id,
  output [7:0]  io_out_aw_bits_len,
  output [2:0]  io_out_aw_bits_size,
  input         io_out_w_ready,
  output        io_out_w_valid,
  output [63:0] io_out_w_bits_data,
  output [7:0]  io_out_w_bits_strb,
  output        io_out_w_bits_last,
  output        io_out_b_ready,
  input         io_out_b_valid,
  input  [3:0]  io_out_b_bits_id,
  input         io_out_ar_ready,
  output        io_out_ar_valid,
  output [31:0] io_out_ar_bits_addr,
  output [3:0]  io_out_ar_bits_id,
  output [7:0]  io_out_ar_bits_len,
  output [2:0]  io_out_ar_bits_size,
  output        io_out_r_ready,
  input         io_out_r_valid,
  input  [63:0] io_out_r_bits_data,
  input  [3:0]  io_out_r_bits_id,
  input         io_out_r_bits_last
);
  wire  _io_out_aw_valid_T = io_in_req_valid & io_in_req_bits_aen; // @[SimpleAxi.scala 48:37]
  wire  _io_in_req_ready_T_1 = io_in_req_bits_wen ? io_out_aw_ready & io_out_w_ready : io_out_ar_ready; // @[SimpleAxi.scala 84:30]
  wire  _io_in_req_ready_T_2 = io_in_req_bits_wen & io_out_w_ready; // @[SimpleAxi.scala 85:30]
  wire [3:0] _io_in_resp_bits_id_T = io_out_r_valid ? io_out_r_bits_id : 4'h0; // @[SimpleAxi.scala 88:28]
  assign io_in_req_ready = io_in_req_bits_aen ? _io_in_req_ready_T_1 : _io_in_req_ready_T_2; // @[SimpleAxi.scala 83:28]
  assign io_in_resp_valid = io_out_b_valid | io_out_r_valid; // @[SimpleAxi.scala 86:37]
  assign io_in_resp_bits_id = io_out_b_valid ? io_out_b_bits_id : _io_in_resp_bits_id_T; // @[SimpleAxi.scala 87:28]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[SimpleAxi.scala 89:22]
  assign io_in_resp_bits_rlast = io_out_r_valid & io_out_r_bits_last; // @[SimpleAxi.scala 91:37]
  assign io_out_aw_valid = io_in_req_valid & io_in_req_bits_aen & io_in_req_bits_wen; // @[SimpleAxi.scala 48:56]
  assign io_out_aw_bits_addr = io_in_req_bits_addr; // @[SimpleAxi.scala 49:21]
  assign io_out_aw_bits_id = io_in_req_bits_id; // @[SimpleAxi.scala 51:21]
  assign io_out_aw_bits_len = io_in_req_bits_len; // @[SimpleAxi.scala 53:21]
  assign io_out_aw_bits_size = {1'h0,io_in_req_bits_size}; // @[Cat.scala 30:58]
  assign io_out_w_valid = io_in_req_valid & io_in_req_bits_wen; // @[SimpleAxi.scala 60:37]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[SimpleAxi.scala 61:21]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[SimpleAxi.scala 62:21]
  assign io_out_w_bits_last = io_in_req_bits_wlast; // @[SimpleAxi.scala 63:21]
  assign io_out_b_ready = io_in_resp_ready; // @[SimpleAxi.scala 79:15]
  assign io_out_ar_valid = _io_out_aw_valid_T & io_in_req_bits_ren; // @[SimpleAxi.scala 65:56]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[SimpleAxi.scala 66:21]
  assign io_out_ar_bits_id = io_in_req_bits_id; // @[SimpleAxi.scala 68:21]
  assign io_out_ar_bits_len = io_in_req_bits_len; // @[SimpleAxi.scala 70:21]
  assign io_out_ar_bits_size = {1'h0,io_in_req_bits_size}; // @[Cat.scala 30:58]
  assign io_out_r_ready = io_in_resp_ready; // @[SimpleAxi.scala 81:15]
endmodule
module ysyx_210340(
  input         clock,
  input         reset,
  input         io_interrupt,
  input         io_master_awready,
  output        io_master_awvalid,
  output [3:0]  io_master_awid,
  output [31:0] io_master_awaddr,
  output [7:0]  io_master_awlen,
  output [2:0]  io_master_awsize,
  output [1:0]  io_master_awburst,
  input         io_master_wready,
  output        io_master_wvalid,
  output [63:0] io_master_wdata,
  output [7:0]  io_master_wstrb,
  output        io_master_wlast,
  output        io_master_bready,
  input         io_master_bvalid,
  input  [3:0]  io_master_bid,
  input  [1:0]  io_master_bresp,
  input         io_master_arready,
  output        io_master_arvalid,
  output [3:0]  io_master_arid,
  output [31:0] io_master_araddr,
  output [7:0]  io_master_arlen,
  output [2:0]  io_master_arsize,
  output [1:0]  io_master_arburst,
  output        io_master_rready,
  input         io_master_rvalid,
  input  [3:0]  io_master_rid,
  input  [1:0]  io_master_rresp,
  input  [63:0] io_master_rdata,
  input         io_master_rlast,
  output        io_slave_awready,
  input         io_slave_awvalid,
  input  [3:0]  io_slave_awid,
  input  [31:0] io_slave_awaddr,
  input  [7:0]  io_slave_awlen,
  input  [2:0]  io_slave_awsize,
  input  [1:0]  io_slave_awburst,
  output        io_slave_wready,
  input         io_slave_wvalid,
  input  [63:0] io_slave_wdata,
  input  [7:0]  io_slave_wstrb,
  input         io_slave_wlast,
  input         io_slave_bready,
  output        io_slave_bvalid,
  output [3:0]  io_slave_bid,
  output [1:0]  io_slave_bresp,
  output        io_slave_arready,
  input         io_slave_arvalid,
  input  [3:0]  io_slave_arid,
  input  [31:0] io_slave_araddr,
  input  [7:0]  io_slave_arlen,
  input  [2:0]  io_slave_arsize,
  input  [1:0]  io_slave_arburst,
  input         io_slave_rready,
  output        io_slave_rvalid,
  output [3:0]  io_slave_rid,
  output [1:0]  io_slave_rresp,
  output [63:0] io_slave_rdata,
  output [5:0]   io_sram0_addr,
  output         io_sram0_cen,
  output         io_sram0_wen,
  output [127:0] io_sram0_wmask,
  output [127:0] io_sram0_wdata,
  input  [127:0] io_sram0_rdata,
  output [5:0]   io_sram1_addr,
  output         io_sram1_cen,
  output         io_sram1_wen,
  output [127:0] io_sram1_wmask,
  output [127:0] io_sram1_wdata,
  input  [127:0] io_sram1_rdata,
  output [5:0]   io_sram2_addr,
  output         io_sram2_cen,
  output         io_sram2_wen,
  output [127:0] io_sram2_wmask,
  output [127:0] io_sram2_wdata,
  input  [127:0] io_sram2_rdata,
  output [5:0]   io_sram3_addr,
  output         io_sram3_cen,
  output         io_sram3_wen,
  output [127:0] io_sram3_wmask,
  output [127:0] io_sram3_wdata,
  input  [127:0] io_sram3_rdata,
  output [5:0]   io_sram4_addr,
  output         io_sram4_cen,
  output         io_sram4_wen,
  output [127:0] io_sram4_wmask,
  output [127:0] io_sram4_wdata,
  input  [127:0] io_sram4_rdata,
  output [5:0]   io_sram5_addr,
  output         io_sram5_cen,
  output         io_sram5_wen,
  output [127:0] io_sram5_wmask,
  output [127:0] io_sram5_wdata,
  input  [127:0] io_sram5_rdata,
  output [5:0]   io_sram6_addr,
  output         io_sram6_cen,
  output         io_sram6_wen,
  output [127:0] io_sram6_wmask,
  output [127:0] io_sram6_wdata,
  input  [127:0] io_sram6_rdata,
  output [5:0]   io_sram7_addr,
  output         io_sram7_cen,
  output         io_sram7_wen,
  output [127:0] io_sram7_wmask,
  output [127:0] io_sram7_wdata,
  input  [127:0] io_sram7_rdata,  
  output        io_slave_rlast
);
  wire  core_clock; // @[SoCTop.scala 13:20]
  wire  core_reset; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_0_req_ready; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_0_req_valid; // @[SoCTop.scala 13:20]
  wire [31:0] core_io_core_bus_0_req_bits_addr; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_0_req_bits_aen; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_0_req_bits_ren; // @[SoCTop.scala 13:20]
  wire [63:0] core_io_core_bus_0_req_bits_wdata; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_0_req_bits_wlast; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_0_req_bits_wen; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_0_resp_ready; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_0_resp_valid; // @[SoCTop.scala 13:20]
  wire [63:0] core_io_core_bus_0_resp_bits_rdata; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_0_resp_bits_rlast; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_1_req_ready; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_1_req_valid; // @[SoCTop.scala 13:20]
  wire [31:0] core_io_core_bus_1_req_bits_addr; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_1_req_bits_aen; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_1_req_bits_ren; // @[SoCTop.scala 13:20]
  wire [63:0] core_io_core_bus_1_req_bits_wdata; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_1_req_bits_wlast; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_1_req_bits_wen; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_1_resp_ready; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_1_resp_valid; // @[SoCTop.scala 13:20]
  wire [63:0] core_io_core_bus_1_resp_bits_rdata; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_1_resp_bits_rlast; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_2_req_ready; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_2_req_valid; // @[SoCTop.scala 13:20]
  wire [31:0] core_io_core_bus_2_req_bits_addr; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_2_req_bits_ren; // @[SoCTop.scala 13:20]
  wire [63:0] core_io_core_bus_2_req_bits_wdata; // @[SoCTop.scala 13:20]
  wire [7:0] core_io_core_bus_2_req_bits_wmask; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_2_req_bits_wen; // @[SoCTop.scala 13:20]
  wire [1:0] core_io_core_bus_2_req_bits_size; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_2_resp_ready; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_2_resp_valid; // @[SoCTop.scala 13:20]
  wire [63:0] core_io_core_bus_2_resp_bits_rdata; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_3_req_ready; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_3_req_valid; // @[SoCTop.scala 13:20]
  wire [31:0] core_io_core_bus_3_req_bits_addr; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_3_req_bits_ren; // @[SoCTop.scala 13:20]
  wire [63:0] core_io_core_bus_3_req_bits_wdata; // @[SoCTop.scala 13:20]
  wire [7:0] core_io_core_bus_3_req_bits_wmask; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_3_req_bits_wen; // @[SoCTop.scala 13:20]
  wire [1:0] core_io_core_bus_3_req_bits_size; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_3_resp_ready; // @[SoCTop.scala 13:20]
  wire  core_io_core_bus_3_resp_valid; // @[SoCTop.scala 13:20]
  wire [63:0] core_io_core_bus_3_resp_bits_rdata; // @[SoCTop.scala 13:20]
  wire  crossbar_clock; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_0_req_ready; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_0_req_valid; // @[SoCTop.scala 15:24]
  wire [31:0] crossbar_io_in_0_req_bits_addr; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_0_req_bits_aen; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_0_req_bits_ren; // @[SoCTop.scala 15:24]
  wire [63:0] crossbar_io_in_0_req_bits_wdata; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_0_req_bits_wlast; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_0_req_bits_wen; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_0_resp_ready; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_0_resp_valid; // @[SoCTop.scala 15:24]
  wire [63:0] crossbar_io_in_0_resp_bits_rdata; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_0_resp_bits_rlast; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_1_req_ready; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_1_req_valid; // @[SoCTop.scala 15:24]
  wire [31:0] crossbar_io_in_1_req_bits_addr; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_1_req_bits_aen; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_1_req_bits_ren; // @[SoCTop.scala 15:24]
  wire [63:0] crossbar_io_in_1_req_bits_wdata; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_1_req_bits_wlast; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_1_req_bits_wen; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_1_resp_ready; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_1_resp_valid; // @[SoCTop.scala 15:24]
  wire [63:0] crossbar_io_in_1_resp_bits_rdata; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_1_resp_bits_rlast; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_2_req_ready; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_2_req_valid; // @[SoCTop.scala 15:24]
  wire [31:0] crossbar_io_in_2_req_bits_addr; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_2_req_bits_ren; // @[SoCTop.scala 15:24]
  wire [63:0] crossbar_io_in_2_req_bits_wdata; // @[SoCTop.scala 15:24]
  wire [7:0] crossbar_io_in_2_req_bits_wmask; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_2_req_bits_wen; // @[SoCTop.scala 15:24]
  wire [1:0] crossbar_io_in_2_req_bits_size; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_2_resp_ready; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_2_resp_valid; // @[SoCTop.scala 15:24]
  wire [63:0] crossbar_io_in_2_resp_bits_rdata; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_3_req_ready; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_3_req_valid; // @[SoCTop.scala 15:24]
  wire [31:0] crossbar_io_in_3_req_bits_addr; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_3_req_bits_ren; // @[SoCTop.scala 15:24]
  wire [63:0] crossbar_io_in_3_req_bits_wdata; // @[SoCTop.scala 15:24]
  wire [7:0] crossbar_io_in_3_req_bits_wmask; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_3_req_bits_wen; // @[SoCTop.scala 15:24]
  wire [1:0] crossbar_io_in_3_req_bits_size; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_3_resp_ready; // @[SoCTop.scala 15:24]
  wire  crossbar_io_in_3_resp_valid; // @[SoCTop.scala 15:24]
  wire [63:0] crossbar_io_in_3_resp_bits_rdata; // @[SoCTop.scala 15:24]
  wire  crossbar_io_out_req_ready; // @[SoCTop.scala 15:24]
  wire  crossbar_io_out_req_valid; // @[SoCTop.scala 15:24]
  wire [3:0] crossbar_io_out_req_bits_id; // @[SoCTop.scala 15:24]
  wire [31:0] crossbar_io_out_req_bits_addr; // @[SoCTop.scala 15:24]
  wire  crossbar_io_out_req_bits_aen; // @[SoCTop.scala 15:24]
  wire  crossbar_io_out_req_bits_ren; // @[SoCTop.scala 15:24]
  wire [63:0] crossbar_io_out_req_bits_wdata; // @[SoCTop.scala 15:24]
  wire [7:0] crossbar_io_out_req_bits_wmask; // @[SoCTop.scala 15:24]
  wire  crossbar_io_out_req_bits_wlast; // @[SoCTop.scala 15:24]
  wire  crossbar_io_out_req_bits_wen; // @[SoCTop.scala 15:24]
  wire [7:0] crossbar_io_out_req_bits_len; // @[SoCTop.scala 15:24]
  wire [1:0] crossbar_io_out_req_bits_size; // @[SoCTop.scala 15:24]
  wire  crossbar_io_out_resp_ready; // @[SoCTop.scala 15:24]
  wire  crossbar_io_out_resp_valid; // @[SoCTop.scala 15:24]
  wire [3:0] crossbar_io_out_resp_bits_id; // @[SoCTop.scala 15:24]
  wire [63:0] crossbar_io_out_resp_bits_rdata; // @[SoCTop.scala 15:24]
  wire  crossbar_io_out_resp_bits_rlast; // @[SoCTop.scala 15:24]
  wire  core2axi_io_in_req_ready; // @[SoCTop.scala 18:24]
  wire  core2axi_io_in_req_valid; // @[SoCTop.scala 18:24]
  wire [3:0] core2axi_io_in_req_bits_id; // @[SoCTop.scala 18:24]
  wire [31:0] core2axi_io_in_req_bits_addr; // @[SoCTop.scala 18:24]
  wire  core2axi_io_in_req_bits_aen; // @[SoCTop.scala 18:24]
  wire  core2axi_io_in_req_bits_ren; // @[SoCTop.scala 18:24]
  wire [63:0] core2axi_io_in_req_bits_wdata; // @[SoCTop.scala 18:24]
  wire [7:0] core2axi_io_in_req_bits_wmask; // @[SoCTop.scala 18:24]
  wire  core2axi_io_in_req_bits_wlast; // @[SoCTop.scala 18:24]
  wire  core2axi_io_in_req_bits_wen; // @[SoCTop.scala 18:24]
  wire [7:0] core2axi_io_in_req_bits_len; // @[SoCTop.scala 18:24]
  wire [1:0] core2axi_io_in_req_bits_size; // @[SoCTop.scala 18:24]
  wire  core2axi_io_in_resp_ready; // @[SoCTop.scala 18:24]
  wire  core2axi_io_in_resp_valid; // @[SoCTop.scala 18:24]
  wire [3:0] core2axi_io_in_resp_bits_id; // @[SoCTop.scala 18:24]
  wire [63:0] core2axi_io_in_resp_bits_rdata; // @[SoCTop.scala 18:24]
  wire  core2axi_io_in_resp_bits_rlast; // @[SoCTop.scala 18:24]
  wire  core2axi_io_out_aw_ready; // @[SoCTop.scala 18:24]
  wire  core2axi_io_out_aw_valid; // @[SoCTop.scala 18:24]
  wire [31:0] core2axi_io_out_aw_bits_addr; // @[SoCTop.scala 18:24]
  wire [3:0] core2axi_io_out_aw_bits_id; // @[SoCTop.scala 18:24]
  wire [7:0] core2axi_io_out_aw_bits_len; // @[SoCTop.scala 18:24]
  wire [2:0] core2axi_io_out_aw_bits_size; // @[SoCTop.scala 18:24]
  wire  core2axi_io_out_w_ready; // @[SoCTop.scala 18:24]
  wire  core2axi_io_out_w_valid; // @[SoCTop.scala 18:24]
  wire [63:0] core2axi_io_out_w_bits_data; // @[SoCTop.scala 18:24]
  wire [7:0] core2axi_io_out_w_bits_strb; // @[SoCTop.scala 18:24]
  wire  core2axi_io_out_w_bits_last; // @[SoCTop.scala 18:24]
  wire  core2axi_io_out_b_ready; // @[SoCTop.scala 18:24]
  wire  core2axi_io_out_b_valid; // @[SoCTop.scala 18:24]
  wire [3:0] core2axi_io_out_b_bits_id; // @[SoCTop.scala 18:24]
  wire  core2axi_io_out_ar_ready; // @[SoCTop.scala 18:24]
  wire  core2axi_io_out_ar_valid; // @[SoCTop.scala 18:24]
  wire [31:0] core2axi_io_out_ar_bits_addr; // @[SoCTop.scala 18:24]
  wire [3:0] core2axi_io_out_ar_bits_id; // @[SoCTop.scala 18:24]
  wire [7:0] core2axi_io_out_ar_bits_len; // @[SoCTop.scala 18:24]
  wire [2:0] core2axi_io_out_ar_bits_size; // @[SoCTop.scala 18:24]
  wire  core2axi_io_out_r_ready; // @[SoCTop.scala 18:24]
  wire  core2axi_io_out_r_valid; // @[SoCTop.scala 18:24]
  wire [63:0] core2axi_io_out_r_bits_data; // @[SoCTop.scala 18:24]
  wire [3:0] core2axi_io_out_r_bits_id; // @[SoCTop.scala 18:24]
  wire  core2axi_io_out_r_bits_last; // @[SoCTop.scala 18:24]

  wire [5:0] icache_io_sram0_addr; 
  wire  icache_io_sram0_cen; 
  wire  icache_io_sram0_wen; 
  wire [127:0] icache_io_sram0_wdata; 
  wire [127:0] icache_io_sram0_rdata; 
  wire [5:0] icache_io_sram1_addr; 
  wire  icache_io_sram1_cen; 
  wire  icache_io_sram1_wen; 
  wire [127:0] icache_io_sram1_wdata; 
  wire [127:0] icache_io_sram1_rdata; 
  wire [5:0] icache_io_sram2_addr; 
  wire  icache_io_sram2_cen; 
  wire  icache_io_sram2_wen; 
  wire [127:0] icache_io_sram2_wdata; 
  wire [127:0] icache_io_sram2_rdata; 
  wire [5:0] icache_io_sram3_addr; 
  wire  icache_io_sram3_cen; 
  wire  icache_io_sram3_wen; 
  wire [127:0] icache_io_sram3_wdata; 
  wire [127:0] icache_io_sram3_rdata; 
  wire [5:0] dcache_io_sram4_addr; 
  wire  dcache_io_sram4_cen; 
  wire  dcache_io_sram4_wen; 
  wire [127:0] dcache_io_sram4_wdata; 
  wire [127:0] dcache_io_sram4_rdata; 
  wire [5:0] dcache_io_sram5_addr; 
  wire  dcache_io_sram5_cen; 
  wire  dcache_io_sram5_wen; 
  wire [127:0] dcache_io_sram5_wdata; 
  wire [127:0] dcache_io_sram5_rdata; 
  wire [5:0] dcache_io_sram6_addr; 
  wire  dcache_io_sram6_cen; 
  wire  dcache_io_sram6_wen; 
  wire [127:0] dcache_io_sram6_wdata; 
  wire [127:0] dcache_io_sram6_rdata; 
  wire [5:0] dcache_io_sram7_addr; 
  wire  dcache_io_sram7_cen; 
  wire  dcache_io_sram7_wen; 
  wire [127:0] dcache_io_sram7_wdata; 
  wire [127:0] dcache_io_sram7_rdata; 

  ysyx_210340_Core core ( // @[SoCTop.scala 13:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_sram0_cen(icache_io_sram0_cen), 
    .io_sram0_wen(icache_io_sram0_wen), 
    .io_sram0_addr(icache_io_sram0_addr), 
    .io_sram0_wdata(icache_io_sram0_wdata), 
    .io_sram0_rdata(icache_io_sram0_rdata), 
    .io_sram1_cen(icache_io_sram1_cen), 
    .io_sram1_wen(icache_io_sram1_wen), 
    .io_sram1_addr(icache_io_sram1_addr), 
    .io_sram1_wdata(icache_io_sram1_wdata), 
    .io_sram1_rdata(icache_io_sram1_rdata),  
    .io_sram2_cen(icache_io_sram2_cen), 
    .io_sram2_wen(icache_io_sram2_wen), 
    .io_sram2_addr(icache_io_sram2_addr), 
    .io_sram2_wdata(icache_io_sram2_wdata), 
    .io_sram2_rdata(icache_io_sram2_rdata),   
    .io_sram3_cen(icache_io_sram3_cen), 
    .io_sram3_wen(icache_io_sram3_wen), 
    .io_sram3_addr(icache_io_sram3_addr), 
    .io_sram3_wdata(icache_io_sram3_wdata), 
    .io_sram3_rdata(icache_io_sram3_rdata),  
    .io_sram4_cen(dcache_io_sram4_cen), 
    .io_sram4_wen(dcache_io_sram4_wen), 
    .io_sram4_addr(dcache_io_sram4_addr), 
    .io_sram4_wdata(dcache_io_sram4_wdata), 
    .io_sram4_rdata(dcache_io_sram4_rdata), 
    .io_sram5_cen(dcache_io_sram5_cen), 
    .io_sram5_wen(dcache_io_sram5_wen), 
    .io_sram5_addr(dcache_io_sram5_addr), 
    .io_sram5_wdata(dcache_io_sram5_wdata), 
    .io_sram5_rdata(dcache_io_sram5_rdata), 
    .io_sram6_cen(dcache_io_sram6_cen), 
    .io_sram6_wen(dcache_io_sram6_wen), 
    .io_sram6_addr(dcache_io_sram6_addr), 
    .io_sram6_wdata(dcache_io_sram6_wdata), 
    .io_sram6_rdata(dcache_io_sram6_rdata),   
    .io_sram7_cen(dcache_io_sram7_cen), 
    .io_sram7_wen(dcache_io_sram7_wen), 
    .io_sram7_addr(dcache_io_sram7_addr), 
    .io_sram7_wdata(dcache_io_sram7_wdata), 
    .io_sram7_rdata(dcache_io_sram7_rdata),
    .io_core_bus_0_req_ready(core_io_core_bus_0_req_ready),
    .io_core_bus_0_req_valid(core_io_core_bus_0_req_valid),
    .io_core_bus_0_req_bits_addr(core_io_core_bus_0_req_bits_addr),
    .io_core_bus_0_req_bits_aen(core_io_core_bus_0_req_bits_aen),
    .io_core_bus_0_req_bits_ren(core_io_core_bus_0_req_bits_ren),
    .io_core_bus_0_req_bits_wdata(core_io_core_bus_0_req_bits_wdata),
    .io_core_bus_0_req_bits_wlast(core_io_core_bus_0_req_bits_wlast),
    .io_core_bus_0_req_bits_wen(core_io_core_bus_0_req_bits_wen),
    .io_core_bus_0_resp_ready(core_io_core_bus_0_resp_ready),
    .io_core_bus_0_resp_valid(core_io_core_bus_0_resp_valid),
    .io_core_bus_0_resp_bits_rdata(core_io_core_bus_0_resp_bits_rdata),
    .io_core_bus_0_resp_bits_rlast(core_io_core_bus_0_resp_bits_rlast),
    .io_core_bus_1_req_ready(core_io_core_bus_1_req_ready),
    .io_core_bus_1_req_valid(core_io_core_bus_1_req_valid),
    .io_core_bus_1_req_bits_addr(core_io_core_bus_1_req_bits_addr),
    .io_core_bus_1_req_bits_aen(core_io_core_bus_1_req_bits_aen),
    .io_core_bus_1_req_bits_ren(core_io_core_bus_1_req_bits_ren),
    .io_core_bus_1_req_bits_wdata(core_io_core_bus_1_req_bits_wdata),
    .io_core_bus_1_req_bits_wlast(core_io_core_bus_1_req_bits_wlast),
    .io_core_bus_1_req_bits_wen(core_io_core_bus_1_req_bits_wen),
    .io_core_bus_1_resp_ready(core_io_core_bus_1_resp_ready),
    .io_core_bus_1_resp_valid(core_io_core_bus_1_resp_valid),
    .io_core_bus_1_resp_bits_rdata(core_io_core_bus_1_resp_bits_rdata),
    .io_core_bus_1_resp_bits_rlast(core_io_core_bus_1_resp_bits_rlast),
    .io_core_bus_2_req_ready(core_io_core_bus_2_req_ready),
    .io_core_bus_2_req_valid(core_io_core_bus_2_req_valid),
    .io_core_bus_2_req_bits_addr(core_io_core_bus_2_req_bits_addr),
    .io_core_bus_2_req_bits_ren(core_io_core_bus_2_req_bits_ren),
    .io_core_bus_2_req_bits_wdata(core_io_core_bus_2_req_bits_wdata),
    .io_core_bus_2_req_bits_wmask(core_io_core_bus_2_req_bits_wmask),
    .io_core_bus_2_req_bits_wen(core_io_core_bus_2_req_bits_wen),
    .io_core_bus_2_req_bits_size(core_io_core_bus_2_req_bits_size),
    .io_core_bus_2_resp_ready(core_io_core_bus_2_resp_ready),
    .io_core_bus_2_resp_valid(core_io_core_bus_2_resp_valid),
    .io_core_bus_2_resp_bits_rdata(core_io_core_bus_2_resp_bits_rdata),
    .io_core_bus_3_req_ready(core_io_core_bus_3_req_ready),
    .io_core_bus_3_req_valid(core_io_core_bus_3_req_valid),
    .io_core_bus_3_req_bits_addr(core_io_core_bus_3_req_bits_addr),
    .io_core_bus_3_req_bits_ren(core_io_core_bus_3_req_bits_ren),
    .io_core_bus_3_req_bits_wdata(core_io_core_bus_3_req_bits_wdata),
    .io_core_bus_3_req_bits_wmask(core_io_core_bus_3_req_bits_wmask),
    .io_core_bus_3_req_bits_wen(core_io_core_bus_3_req_bits_wen),
    .io_core_bus_3_req_bits_size(core_io_core_bus_3_req_bits_size),
    .io_core_bus_3_resp_ready(core_io_core_bus_3_resp_ready),
    .io_core_bus_3_resp_valid(core_io_core_bus_3_resp_valid),
    .io_core_bus_3_resp_bits_rdata(core_io_core_bus_3_resp_bits_rdata)
  );

  assign io_sram0_wmask = 128'h0000000000000000;
  assign io_sram1_wmask = 128'h0000000000000000;
  assign io_sram2_wmask = 128'h0000000000000000;
  assign io_sram3_wmask = 128'h0000000000000000;
  assign io_sram4_wmask = 128'h0000000000000000;
  assign io_sram5_wmask = 128'h0000000000000000;
  assign io_sram6_wmask = 128'h0000000000000000;
  assign io_sram7_wmask = 128'h0000000000000000;

  assign io_sram0_addr = icache_io_sram0_addr; // @[cpu.scala 163:22]
  assign io_sram0_cen = icache_io_sram0_cen; // @[cpu.scala 163:22]
  assign io_sram0_wen = icache_io_sram0_wen; // @[cpu.scala 163:22]
  assign io_sram0_wdata = icache_io_sram0_wdata; // @[cpu.scala 163:22]
  assign io_sram1_addr = icache_io_sram1_addr; // @[cpu.scala 164:22]
  assign io_sram1_cen = icache_io_sram1_cen; // @[cpu.scala 164:22]
  assign io_sram1_wen = icache_io_sram1_wen; // @[cpu.scala 164:22]
  assign io_sram1_wdata = icache_io_sram1_wdata; // @[cpu.scala 164:22]
  assign io_sram2_addr = icache_io_sram2_addr; // @[cpu.scala 165:22]
  assign io_sram2_cen = icache_io_sram2_cen; // @[cpu.scala 165:22]
  assign io_sram2_wen = icache_io_sram2_wen; // @[cpu.scala 165:22]
  assign io_sram2_wdata = icache_io_sram2_wdata; // @[cpu.scala 165:22]
  assign io_sram3_addr = icache_io_sram3_addr; // @[cpu.scala 166:22]
  assign io_sram3_cen = icache_io_sram3_cen; // @[cpu.scala 166:22]
  assign io_sram3_wen = icache_io_sram3_wen; // @[cpu.scala 166:22]
  assign io_sram3_wdata = icache_io_sram3_wdata; // @[cpu.scala 166:22]
  assign io_sram4_addr = dcache_io_sram4_addr; // @[cpu.scala 167:22]
  assign io_sram4_cen = dcache_io_sram4_cen; // @[cpu.scala 167:22]
  assign io_sram4_wen = dcache_io_sram4_wen; // @[cpu.scala 167:22]
  assign io_sram4_wdata = dcache_io_sram4_wdata; // @[cpu.scala 167:22]
  assign io_sram5_addr = dcache_io_sram5_addr; // @[cpu.scala 168:22]
  assign io_sram5_cen = dcache_io_sram5_cen; // @[cpu.scala 168:22]
  assign io_sram5_wen = dcache_io_sram5_wen; // @[cpu.scala 168:22]
  assign io_sram5_wdata = dcache_io_sram5_wdata; // @[cpu.scala 168:22]
  assign io_sram6_addr = dcache_io_sram6_addr; // @[cpu.scala 169:22]
  assign io_sram6_cen = dcache_io_sram6_cen; // @[cpu.scala 169:22]
  assign io_sram6_wen = dcache_io_sram6_wen; // @[cpu.scala 169:22]
  assign io_sram6_wdata = dcache_io_sram6_wdata; // @[cpu.scala 169:22]
  assign io_sram7_addr = dcache_io_sram7_addr; // @[cpu.scala 170:22]
  assign io_sram7_cen = dcache_io_sram7_cen; // @[cpu.scala 170:22]
  assign io_sram7_wen = dcache_io_sram7_wen; // @[cpu.scala 170:22]
  assign io_sram7_wdata = dcache_io_sram7_wdata; // @[cpu.scala 170:22]

  assign icache_io_sram0_rdata = io_sram0_rdata;
  assign icache_io_sram1_rdata = io_sram1_rdata;
  assign icache_io_sram2_rdata = io_sram2_rdata;
  assign icache_io_sram3_rdata = io_sram3_rdata;
  assign dcache_io_sram4_rdata = io_sram4_rdata;
  assign dcache_io_sram5_rdata = io_sram5_rdata;
  assign dcache_io_sram6_rdata = io_sram6_rdata;
  assign dcache_io_sram7_rdata = io_sram7_rdata;

  ysyx_210340_CoreBusCrossbarNto1 crossbar ( // @[SoCTop.scala 15:24]
    .clock(crossbar_clock),
    .io_in_0_req_ready(crossbar_io_in_0_req_ready),
    .io_in_0_req_valid(crossbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(crossbar_io_in_0_req_bits_addr),
    .io_in_0_req_bits_aen(crossbar_io_in_0_req_bits_aen),
    .io_in_0_req_bits_ren(crossbar_io_in_0_req_bits_ren),
    .io_in_0_req_bits_wdata(crossbar_io_in_0_req_bits_wdata),
    .io_in_0_req_bits_wlast(crossbar_io_in_0_req_bits_wlast),
    .io_in_0_req_bits_wen(crossbar_io_in_0_req_bits_wen),
    .io_in_0_resp_ready(crossbar_io_in_0_resp_ready),
    .io_in_0_resp_valid(crossbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_rdata(crossbar_io_in_0_resp_bits_rdata),
    .io_in_0_resp_bits_rlast(crossbar_io_in_0_resp_bits_rlast),
    .io_in_1_req_ready(crossbar_io_in_1_req_ready),
    .io_in_1_req_valid(crossbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(crossbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_aen(crossbar_io_in_1_req_bits_aen),
    .io_in_1_req_bits_ren(crossbar_io_in_1_req_bits_ren),
    .io_in_1_req_bits_wdata(crossbar_io_in_1_req_bits_wdata),
    .io_in_1_req_bits_wlast(crossbar_io_in_1_req_bits_wlast),
    .io_in_1_req_bits_wen(crossbar_io_in_1_req_bits_wen),
    .io_in_1_resp_ready(crossbar_io_in_1_resp_ready),
    .io_in_1_resp_valid(crossbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_rdata(crossbar_io_in_1_resp_bits_rdata),
    .io_in_1_resp_bits_rlast(crossbar_io_in_1_resp_bits_rlast),
    .io_in_2_req_ready(crossbar_io_in_2_req_ready),
    .io_in_2_req_valid(crossbar_io_in_2_req_valid),
    .io_in_2_req_bits_addr(crossbar_io_in_2_req_bits_addr),
    .io_in_2_req_bits_ren(crossbar_io_in_2_req_bits_ren),
    .io_in_2_req_bits_wdata(crossbar_io_in_2_req_bits_wdata),
    .io_in_2_req_bits_wmask(crossbar_io_in_2_req_bits_wmask),
    .io_in_2_req_bits_wen(crossbar_io_in_2_req_bits_wen),
    .io_in_2_req_bits_size(crossbar_io_in_2_req_bits_size),
    .io_in_2_resp_ready(crossbar_io_in_2_resp_ready),
    .io_in_2_resp_valid(crossbar_io_in_2_resp_valid),
    .io_in_2_resp_bits_rdata(crossbar_io_in_2_resp_bits_rdata),
    .io_in_3_req_ready(crossbar_io_in_3_req_ready),
    .io_in_3_req_valid(crossbar_io_in_3_req_valid),
    .io_in_3_req_bits_addr(crossbar_io_in_3_req_bits_addr),
    .io_in_3_req_bits_ren(crossbar_io_in_3_req_bits_ren),
    .io_in_3_req_bits_wdata(crossbar_io_in_3_req_bits_wdata),
    .io_in_3_req_bits_wmask(crossbar_io_in_3_req_bits_wmask),
    .io_in_3_req_bits_wen(crossbar_io_in_3_req_bits_wen),
    .io_in_3_req_bits_size(crossbar_io_in_3_req_bits_size),
    .io_in_3_resp_ready(crossbar_io_in_3_resp_ready),
    .io_in_3_resp_valid(crossbar_io_in_3_resp_valid),
    .io_in_3_resp_bits_rdata(crossbar_io_in_3_resp_bits_rdata),
    .io_out_req_ready(crossbar_io_out_req_ready),
    .io_out_req_valid(crossbar_io_out_req_valid),
    .io_out_req_bits_id(crossbar_io_out_req_bits_id),
    .io_out_req_bits_addr(crossbar_io_out_req_bits_addr),
    .io_out_req_bits_aen(crossbar_io_out_req_bits_aen),
    .io_out_req_bits_ren(crossbar_io_out_req_bits_ren),
    .io_out_req_bits_wdata(crossbar_io_out_req_bits_wdata),
    .io_out_req_bits_wmask(crossbar_io_out_req_bits_wmask),
    .io_out_req_bits_wlast(crossbar_io_out_req_bits_wlast),
    .io_out_req_bits_wen(crossbar_io_out_req_bits_wen),
    .io_out_req_bits_len(crossbar_io_out_req_bits_len),
    .io_out_req_bits_size(crossbar_io_out_req_bits_size),
    .io_out_resp_ready(crossbar_io_out_resp_ready),
    .io_out_resp_valid(crossbar_io_out_resp_valid),
    .io_out_resp_bits_id(crossbar_io_out_resp_bits_id),
    .io_out_resp_bits_rdata(crossbar_io_out_resp_bits_rdata),
    .io_out_resp_bits_rlast(crossbar_io_out_resp_bits_rlast)
  );
  ysyx_210340_SimpleAxi2Axi core2axi ( // @[SoCTop.scala 18:24]
    .io_in_req_ready(core2axi_io_in_req_ready),
    .io_in_req_valid(core2axi_io_in_req_valid),
    .io_in_req_bits_id(core2axi_io_in_req_bits_id),
    .io_in_req_bits_addr(core2axi_io_in_req_bits_addr),
    .io_in_req_bits_aen(core2axi_io_in_req_bits_aen),
    .io_in_req_bits_ren(core2axi_io_in_req_bits_ren),
    .io_in_req_bits_wdata(core2axi_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(core2axi_io_in_req_bits_wmask),
    .io_in_req_bits_wlast(core2axi_io_in_req_bits_wlast),
    .io_in_req_bits_wen(core2axi_io_in_req_bits_wen),
    .io_in_req_bits_len(core2axi_io_in_req_bits_len),
    .io_in_req_bits_size(core2axi_io_in_req_bits_size),
    .io_in_resp_ready(core2axi_io_in_resp_ready),
    .io_in_resp_valid(core2axi_io_in_resp_valid),
    .io_in_resp_bits_id(core2axi_io_in_resp_bits_id),
    .io_in_resp_bits_rdata(core2axi_io_in_resp_bits_rdata),
    .io_in_resp_bits_rlast(core2axi_io_in_resp_bits_rlast),
    .io_out_aw_ready(core2axi_io_out_aw_ready),
    .io_out_aw_valid(core2axi_io_out_aw_valid),
    .io_out_aw_bits_addr(core2axi_io_out_aw_bits_addr),
    .io_out_aw_bits_id(core2axi_io_out_aw_bits_id),
    .io_out_aw_bits_len(core2axi_io_out_aw_bits_len),
    .io_out_aw_bits_size(core2axi_io_out_aw_bits_size),
    .io_out_w_ready(core2axi_io_out_w_ready),
    .io_out_w_valid(core2axi_io_out_w_valid),
    .io_out_w_bits_data(core2axi_io_out_w_bits_data),
    .io_out_w_bits_strb(core2axi_io_out_w_bits_strb),
    .io_out_w_bits_last(core2axi_io_out_w_bits_last),
    .io_out_b_ready(core2axi_io_out_b_ready),
    .io_out_b_valid(core2axi_io_out_b_valid),
    .io_out_b_bits_id(core2axi_io_out_b_bits_id),
    .io_out_ar_ready(core2axi_io_out_ar_ready),
    .io_out_ar_valid(core2axi_io_out_ar_valid),
    .io_out_ar_bits_addr(core2axi_io_out_ar_bits_addr),
    .io_out_ar_bits_id(core2axi_io_out_ar_bits_id),
    .io_out_ar_bits_len(core2axi_io_out_ar_bits_len),
    .io_out_ar_bits_size(core2axi_io_out_ar_bits_size),
    .io_out_r_ready(core2axi_io_out_r_ready),
    .io_out_r_valid(core2axi_io_out_r_valid),
    .io_out_r_bits_data(core2axi_io_out_r_bits_data),
    .io_out_r_bits_id(core2axi_io_out_r_bits_id),
    .io_out_r_bits_last(core2axi_io_out_r_bits_last)
  );
  assign io_master_awvalid = core2axi_io_out_aw_valid; // @[SoCTop.scala 20:16]
  assign io_master_awid = core2axi_io_out_aw_bits_id; // @[SoCTop.scala 20:16]
  assign io_master_awaddr = core2axi_io_out_aw_bits_addr; // @[SoCTop.scala 20:16]
  assign io_master_awlen = core2axi_io_out_aw_bits_len; // @[SoCTop.scala 20:16]
  assign io_master_awsize = core2axi_io_out_aw_bits_size; // @[SoCTop.scala 20:16]
  assign io_master_awburst = 2'h1; // @[SoCTop.scala 20:16]
  assign io_master_wvalid = core2axi_io_out_w_valid; // @[SoCTop.scala 20:16]
  assign io_master_wdata = core2axi_io_out_w_bits_data; // @[SoCTop.scala 20:16]
  assign io_master_wstrb = core2axi_io_out_w_bits_strb; // @[SoCTop.scala 20:16]
  assign io_master_wlast = core2axi_io_out_w_bits_last; // @[SoCTop.scala 20:16]
  assign io_master_bready = core2axi_io_out_b_ready; // @[SoCTop.scala 20:16]
  assign io_master_arvalid = core2axi_io_out_ar_valid; // @[SoCTop.scala 20:16]
  assign io_master_arid = core2axi_io_out_ar_bits_id; // @[SoCTop.scala 20:16]
  assign io_master_araddr = core2axi_io_out_ar_bits_addr; // @[SoCTop.scala 20:16]
  assign io_master_arlen = core2axi_io_out_ar_bits_len; // @[SoCTop.scala 20:16]
  assign io_master_arsize = core2axi_io_out_ar_bits_size; // @[SoCTop.scala 20:16]
  assign io_master_arburst = 2'h1; // @[SoCTop.scala 20:16]
  assign io_master_rready = core2axi_io_out_r_ready; // @[SoCTop.scala 20:16]
  assign io_slave_awready = 1'h0; // @[SoCTop.scala 23:21]
  assign io_slave_wready = 1'h0; // @[SoCTop.scala 24:21]
  assign io_slave_bvalid = 1'h0; // @[SoCTop.scala 25:21]
  assign io_slave_bid = 4'h0; // @[SoCTop.scala 27:21]
  assign io_slave_bresp = 2'h0; // @[SoCTop.scala 26:21]
  assign io_slave_arready = 1'h0; // @[SoCTop.scala 28:21]
  assign io_slave_rvalid = 1'h0; // @[SoCTop.scala 29:21]
  assign io_slave_rid = 4'h0; // @[SoCTop.scala 33:21]
  assign io_slave_rresp = 2'h0; // @[SoCTop.scala 30:21]
  assign io_slave_rdata = 64'h0; // @[SoCTop.scala 31:21]
  assign io_slave_rlast = 1'h0; // @[SoCTop.scala 32:21]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_core_bus_0_req_ready = crossbar_io_in_0_req_ready; // @[SoCTop.scala 16:18]
  assign core_io_core_bus_0_resp_valid = crossbar_io_in_0_resp_valid; // @[SoCTop.scala 16:18]
  assign core_io_core_bus_0_resp_bits_rdata = crossbar_io_in_0_resp_bits_rdata; // @[SoCTop.scala 16:18]
  assign core_io_core_bus_0_resp_bits_rlast = crossbar_io_in_0_resp_bits_rlast; // @[SoCTop.scala 16:18]
  assign core_io_core_bus_1_req_ready = crossbar_io_in_1_req_ready; // @[SoCTop.scala 16:18]
  assign core_io_core_bus_1_resp_valid = crossbar_io_in_1_resp_valid; // @[SoCTop.scala 16:18]
  assign core_io_core_bus_1_resp_bits_rdata = crossbar_io_in_1_resp_bits_rdata; // @[SoCTop.scala 16:18]
  assign core_io_core_bus_1_resp_bits_rlast = crossbar_io_in_1_resp_bits_rlast; // @[SoCTop.scala 16:18]
  assign core_io_core_bus_2_req_ready = crossbar_io_in_2_req_ready; // @[SoCTop.scala 16:18]
  assign core_io_core_bus_2_resp_valid = crossbar_io_in_2_resp_valid; // @[SoCTop.scala 16:18]
  assign core_io_core_bus_2_resp_bits_rdata = crossbar_io_in_2_resp_bits_rdata; // @[SoCTop.scala 16:18]
  assign core_io_core_bus_3_req_ready = crossbar_io_in_3_req_ready; // @[SoCTop.scala 16:18]
  assign core_io_core_bus_3_resp_valid = crossbar_io_in_3_resp_valid; // @[SoCTop.scala 16:18]
  assign core_io_core_bus_3_resp_bits_rdata = crossbar_io_in_3_resp_bits_rdata; // @[SoCTop.scala 16:18]
  assign crossbar_clock = clock;
  assign crossbar_io_in_0_req_valid = core_io_core_bus_0_req_valid; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_0_req_bits_addr = core_io_core_bus_0_req_bits_addr; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_0_req_bits_aen = core_io_core_bus_0_req_bits_aen; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_0_req_bits_ren = core_io_core_bus_0_req_bits_ren; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_0_req_bits_wdata = core_io_core_bus_0_req_bits_wdata; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_0_req_bits_wlast = core_io_core_bus_0_req_bits_wlast; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_0_req_bits_wen = core_io_core_bus_0_req_bits_wen; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_0_resp_ready = core_io_core_bus_0_resp_ready; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_1_req_valid = core_io_core_bus_1_req_valid; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_1_req_bits_addr = core_io_core_bus_1_req_bits_addr; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_1_req_bits_aen = core_io_core_bus_1_req_bits_aen; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_1_req_bits_ren = core_io_core_bus_1_req_bits_ren; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_1_req_bits_wdata = core_io_core_bus_1_req_bits_wdata; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_1_req_bits_wlast = core_io_core_bus_1_req_bits_wlast; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_1_req_bits_wen = core_io_core_bus_1_req_bits_wen; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_1_resp_ready = core_io_core_bus_1_resp_ready; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_2_req_valid = core_io_core_bus_2_req_valid; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_2_req_bits_addr = core_io_core_bus_2_req_bits_addr; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_2_req_bits_ren = core_io_core_bus_2_req_bits_ren; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_2_req_bits_wdata = core_io_core_bus_2_req_bits_wdata; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_2_req_bits_wmask = core_io_core_bus_2_req_bits_wmask; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_2_req_bits_wen = core_io_core_bus_2_req_bits_wen; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_2_req_bits_size = core_io_core_bus_2_req_bits_size; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_2_resp_ready = core_io_core_bus_2_resp_ready; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_3_req_valid = core_io_core_bus_3_req_valid; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_3_req_bits_addr = core_io_core_bus_3_req_bits_addr; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_3_req_bits_ren = core_io_core_bus_3_req_bits_ren; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_3_req_bits_wdata = core_io_core_bus_3_req_bits_wdata; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_3_req_bits_wmask = core_io_core_bus_3_req_bits_wmask; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_3_req_bits_wen = core_io_core_bus_3_req_bits_wen; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_3_req_bits_size = core_io_core_bus_3_req_bits_size; // @[SoCTop.scala 16:18]
  assign crossbar_io_in_3_resp_ready = core_io_core_bus_3_resp_ready; // @[SoCTop.scala 16:18]
  assign crossbar_io_out_req_ready = core2axi_io_in_req_ready; // @[SoCTop.scala 19:15]
  assign crossbar_io_out_resp_valid = core2axi_io_in_resp_valid; // @[SoCTop.scala 19:15]
  assign crossbar_io_out_resp_bits_id = core2axi_io_in_resp_bits_id; // @[SoCTop.scala 19:15]
  assign crossbar_io_out_resp_bits_rdata = core2axi_io_in_resp_bits_rdata; // @[SoCTop.scala 19:15]
  assign crossbar_io_out_resp_bits_rlast = core2axi_io_in_resp_bits_rlast; // @[SoCTop.scala 19:15]
  assign core2axi_io_in_req_valid = crossbar_io_out_req_valid; // @[SoCTop.scala 19:15]
  assign core2axi_io_in_req_bits_id = crossbar_io_out_req_bits_id; // @[SoCTop.scala 19:15]
  assign core2axi_io_in_req_bits_addr = crossbar_io_out_req_bits_addr; // @[SoCTop.scala 19:15]
  assign core2axi_io_in_req_bits_aen = crossbar_io_out_req_bits_aen; // @[SoCTop.scala 19:15]
  assign core2axi_io_in_req_bits_ren = crossbar_io_out_req_bits_ren; // @[SoCTop.scala 19:15]
  assign core2axi_io_in_req_bits_wdata = crossbar_io_out_req_bits_wdata; // @[SoCTop.scala 19:15]
  assign core2axi_io_in_req_bits_wmask = crossbar_io_out_req_bits_wmask; // @[SoCTop.scala 19:15]
  assign core2axi_io_in_req_bits_wlast = crossbar_io_out_req_bits_wlast; // @[SoCTop.scala 19:15]
  assign core2axi_io_in_req_bits_wen = crossbar_io_out_req_bits_wen; // @[SoCTop.scala 19:15]
  assign core2axi_io_in_req_bits_len = crossbar_io_out_req_bits_len; // @[SoCTop.scala 19:15]
  assign core2axi_io_in_req_bits_size = crossbar_io_out_req_bits_size; // @[SoCTop.scala 19:15]
  assign core2axi_io_in_resp_ready = crossbar_io_out_resp_ready; // @[SoCTop.scala 19:15]
  assign core2axi_io_out_aw_ready = io_master_awready; // @[SoCTop.scala 20:16]
  assign core2axi_io_out_w_ready = io_master_wready; // @[SoCTop.scala 20:16]
  assign core2axi_io_out_b_valid = io_master_bvalid; // @[SoCTop.scala 20:16]
  assign core2axi_io_out_b_bits_id = io_master_bid; // @[SoCTop.scala 20:16]
  assign core2axi_io_out_ar_ready = io_master_arready; // @[SoCTop.scala 20:16]
  assign core2axi_io_out_r_valid = io_master_rvalid; // @[SoCTop.scala 20:16]
  assign core2axi_io_out_r_bits_data = io_master_rdata; // @[SoCTop.scala 20:16]
  assign core2axi_io_out_r_bits_id = io_master_rid; // @[SoCTop.scala 20:16]
  assign core2axi_io_out_r_bits_last = io_master_rlast; // @[SoCTop.scala 20:16]
endmodule
