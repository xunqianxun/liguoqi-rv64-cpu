module ysyx_210539_Fetch(
  input         clock,
  input         reset,
  output [31:0] io_instRead_addr,
  input  [63:0] io_instRead_inst,
  output        io_instRead_arvalid,
  input         io_instRead_rvalid,
  output [63:0] io_va2pa_vaddr,
  output        io_va2pa_vvalid,
  input  [31:0] io_va2pa_paddr,
  input         io_va2pa_pvalid,
  input  [63:0] io_va2pa_tlb_excep_cause,
  input  [63:0] io_va2pa_tlb_excep_tval,
  input         io_va2pa_tlb_excep_en,
  input  [63:0] io_reg2if_seq_pc,
  input         io_reg2if_valid,
  input  [63:0] io_wb2if_seq_pc,
  input         io_wb2if_valid,
  input         io_recov,
  input         io_intr_in_en,
  input  [63:0] io_intr_in_cause,
  input  [63:0] io_branchFail_seq_pc,
  input         io_branchFail_valid,
  output [31:0] io_if2id_inst,
  output [63:0] io_if2id_pc,
  output [63:0] io_if2id_excep_cause,
  output [63:0] io_if2id_excep_tval,
  output        io_if2id_excep_en,
  output [63:0] io_if2id_excep_pc,
  input         io_if2id_drop,
  input         io_if2id_stall,
  output        io_if2id_recov,
  output        io_if2id_valid,
  input         io_if2id_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [127:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] pc; // @[fetch.scala 61:21]
  reg  drop1_r; // @[fetch.scala 63:26]
  reg  drop2_r; // @[fetch.scala 64:26]
  reg  drop3_r; // @[fetch.scala 65:26]
  reg  stall1_r; // @[fetch.scala 66:27]
  reg  stall2_r; // @[fetch.scala 67:27]
  reg  stall3_r; // @[fetch.scala 68:27]
  reg  recov3_r; // @[fetch.scala 71:27]
  wire  drop3_in = drop3_r | io_if2id_drop; // @[fetch.scala 83:28]
  wire  drop2_in = drop2_r | drop3_in; // @[fetch.scala 84:28]
  wire  drop1_in = drop1_r | drop2_in; // @[fetch.scala 85:28]
  wire  _stall3_in_T = ~io_if2id_drop; // @[fetch.scala 86:34]
  wire  stall3_in = stall3_r & ~io_if2id_drop | io_if2id_stall; // @[fetch.scala 86:50]
  wire  _stall2_in_T = ~drop3_in; // @[fetch.scala 87:34]
  wire  stall2_in = stall2_r & ~drop3_in | stall3_in; // @[fetch.scala 87:45]
  wire  _stall1_in_T = ~drop2_in; // @[fetch.scala 88:34]
  wire  stall1_in = stall1_r & ~drop2_in | stall2_in; // @[fetch.scala 88:45]
  reg  state; // @[fetch.scala 91:24]
  wire  _T = ~state; // @[Conditional.scala 37:30]
  wire  _GEN_0 = stall1_in | state; // @[fetch.scala 94:28 fetch.scala 95:23 fetch.scala 91:24]
  reg [63:0] pc1_r; // @[fetch.scala 105:24]
  reg [63:0] excep1_r_cause; // @[fetch.scala 107:30]
  reg  excep1_r_en; // @[fetch.scala 107:30]
  reg  valid1_r; // @[fetch.scala 108:30]
  wire  hs_in = _T & ~drop1_in; // @[fetch.scala 109:39]
  wire [63:0] _cur_pc_T_1 = pc + 64'h8; // @[fetch.scala 114:40]
  reg  valid2_r; // @[fetch.scala 156:30]
  reg [1:0] buf_bitmap; // @[fetch.scala 212:34]
  wire  _T_14 = buf_bitmap == 2'h3; // @[fetch.scala 228:25]
  reg  excep_buf_en; // @[fetch.scala 213:34]
  reg  excep2_r_en; // @[fetch.scala 157:30]
  reg  reset_ic; // @[fetch.scala 217:30]
  wire  _T_19 = valid2_r & io_instRead_rvalid & ~reset_ic; // @[fetch.scala 233:51]
  wire  _GEN_76 = excep2_r_en & valid2_r | _T_19; // @[fetch.scala 229:44 fetch.scala 231:17]
  wire  _GEN_88 = buf_bitmap == 2'h3 | excep_buf_en ? 1'h0 : _GEN_76; // @[fetch.scala 228:49 fetch.scala 222:9]
  wire  hs2 = _stall2_in_T & _GEN_88; // @[fetch.scala 227:20 fetch.scala 222:9]
  reg  reset_tlb; // @[fetch.scala 161:30]
  wire  _tlb_inp_valid_T_1 = io_va2pa_pvalid | io_va2pa_tlb_excep_en; // @[fetch.scala 166:58]
  wire  tlb_inp_valid = ~reset_tlb & (io_va2pa_pvalid | io_va2pa_tlb_excep_en); // @[fetch.scala 166:38]
  wire  _GEN_16 = (tlb_inp_valid | excep1_r_en) & valid1_r; // @[fetch.scala 172:49 fetch.scala 173:17 fetch.scala 168:9]
  wire  _GEN_17 = valid2_r & ~hs2 ? 1'h0 : _GEN_16; // @[fetch.scala 170:31 fetch.scala 171:17]
  wire  hs1 = _stall1_in_T & _GEN_17; // @[fetch.scala 169:20 fetch.scala 168:9]
  wire [63:0] cur_pc = hs1 ? _cur_pc_T_1 : pc; // @[Mux.scala 47:69]
  wire [63:0] _next_pc_T = io_branchFail_valid ? io_branchFail_seq_pc : cur_pc; // @[Mux.scala 47:69]
  wire  _GEN_10 = hs_in & io_intr_in_en; // @[fetch.scala 126:16 fetch.scala 72:13]
  wire  _GEN_12 = hs1 ? 1'h0 : valid1_r; // @[fetch.scala 141:24 fetch.scala 142:22 fetch.scala 108:30]
  wire  _GEN_13 = hs_in | _GEN_12; // @[fetch.scala 139:20 fetch.scala 140:22]
  wire  _GEN_14 = _stall1_in_T & _GEN_13; // @[fetch.scala 138:20 fetch.scala 145:18]
  reg [63:0] pc2_r; // @[fetch.scala 154:30]
  reg [31:0] paddr2_r; // @[fetch.scala 155:30]
  reg [63:0] excep2_r_cause; // @[fetch.scala 157:30]
  reg [63:0] excep2_r_tval; // @[fetch.scala 157:30]
  reg [63:0] excep2_r_pc; // @[fetch.scala 157:30]
  wire  _GEN_19 = hs2 ? 1'h0 : valid2_r; // @[fetch.scala 181:24 fetch.scala 182:22 fetch.scala 156:30]
  wire  _GEN_20 = hs1 | _GEN_19; // @[fetch.scala 177:18 fetch.scala 178:29]
  wire [63:0] _GEN_23 = io_va2pa_tlb_excep_en ? pc1_r : 64'h0; // @[fetch.scala 188:42 fetch.scala 189:28 fetch.scala 195:25]
  wire  _GEN_24 = io_va2pa_tlb_excep_en | excep1_r_en; // @[fetch.scala 188:42 fetch.scala 190:28 fetch.scala 195:25]
  wire [63:0] _GEN_25 = io_va2pa_tlb_excep_en ? io_va2pa_tlb_excep_tval : 64'h0; // @[fetch.scala 188:42 fetch.scala 191:28 fetch.scala 195:25]
  wire [63:0] _GEN_26 = io_va2pa_tlb_excep_en ? io_va2pa_tlb_excep_cause : excep1_r_cause; // @[fetch.scala 188:42 fetch.scala 192:28 fetch.scala 195:25]
  wire  _GEN_35 = io_va2pa_pvalid ? 1'h0 : io_va2pa_tlb_excep_en; // @[fetch.scala 185:36 fetch.scala 72:33]
  wire  _GEN_43 = ~hs1 ? 1'h0 : _GEN_35; // @[fetch.scala 184:19 fetch.scala 72:33]
  wire  _GEN_46 = _stall2_in_T & _GEN_20; // @[fetch.scala 176:20 fetch.scala 198:18]
  wire  _GEN_54 = _stall2_in_T & _GEN_43; // @[fetch.scala 176:20 fetch.scala 72:33]
  wire  cur_excep_en = hs1 ? _GEN_24 : excep2_r_en; // @[fetch.scala 202:27]
  reg [63:0] pc3_r; // @[fetch.scala 205:34]
  reg  valid3_r; // @[fetch.scala 206:34]
  reg [63:0] excep3_r_cause; // @[fetch.scala 207:34]
  reg [63:0] excep3_r_tval; // @[fetch.scala 207:34]
  reg  excep3_r_en; // @[fetch.scala 207:34]
  reg [63:0] excep3_r_pc; // @[fetch.scala 207:34]
  reg [63:0] next_pc_r; // @[fetch.scala 208:34]
  reg  wait_jmp_pc; // @[fetch.scala 209:34]
  reg [127:0] inst_buf; // @[fetch.scala 210:34]
  reg [63:0] buf_start_pc; // @[fetch.scala 211:34]
  reg [63:0] excep_buf_cause; // @[fetch.scala 213:34]
  reg [63:0] excep_buf_tval; // @[fetch.scala 213:34]
  reg [63:0] excep_buf_pc; // @[fetch.scala 213:34]
  reg [31:0] inst_r; // @[fetch.scala 214:34]
  reg  update_excep_pc; // @[fetch.scala 218:34]
  wire [63:0] buf_offset = next_pc_r - buf_start_pc; // @[fetch.scala 223:33]
  wire  hs_out = io_if2id_ready & io_if2id_valid; // @[fetch.scala 224:33]
  wire [63:0] next_inst_buf_lo = inst_buf[63:0]; // @[fetch.scala 236:64]
  wire [127:0] _next_inst_buf_T = {io_instRead_inst,next_inst_buf_lo}; // @[Cat.scala 30:58]
  wire [127:0] _next_inst_buf_T_1 = {64'h0,io_instRead_inst}; // @[Cat.scala 30:58]
  wire [60:0] buf_start_pc_hi = pc2_r[63:3]; // @[fetch.scala 241:42]
  wire [63:0] _buf_start_pc_T = {buf_start_pc_hi,3'h0}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_58 = wait_jmp_pc ? pc2_r : next_pc_r; // @[fetch.scala 242:34 fetch.scala 243:33 fetch.scala 208:34]
  wire  _GEN_59 = wait_jmp_pc ? 1'h0 : wait_jmp_pc; // @[fetch.scala 242:34 fetch.scala 244:33 fetch.scala 209:34]
  wire [127:0] _GEN_60 = buf_bitmap[0] ? _next_inst_buf_T : _next_inst_buf_T_1; // @[fetch.scala 235:32 fetch.scala 236:31 fetch.scala 239:31]
  wire [1:0] _GEN_61 = buf_bitmap[0] ? 2'h3 : 2'h1; // @[fetch.scala 235:32 fetch.scala 237:33 fetch.scala 240:33]
  wire [63:0] _GEN_62 = buf_bitmap[0] ? buf_start_pc : _buf_start_pc_T; // @[fetch.scala 235:32 fetch.scala 211:34 fetch.scala 241:30]
  wire [63:0] _GEN_63 = buf_bitmap[0] ? next_pc_r : _GEN_58; // @[fetch.scala 235:32 fetch.scala 208:34]
  wire  _GEN_64 = buf_bitmap[0] ? wait_jmp_pc : _GEN_59; // @[fetch.scala 235:32 fetch.scala 209:34]
  wire [127:0] _GEN_66 = valid2_r & io_instRead_rvalid & ~reset_ic ? _GEN_60 : inst_buf; // @[fetch.scala 233:64 fetch.scala 225:19]
  wire [1:0] _GEN_67 = valid2_r & io_instRead_rvalid & ~reset_ic ? _GEN_61 : buf_bitmap; // @[fetch.scala 233:64 fetch.scala 226:21]
  wire [63:0] _GEN_68 = valid2_r & io_instRead_rvalid & ~reset_ic ? _GEN_62 : buf_start_pc; // @[fetch.scala 233:64 fetch.scala 211:34]
  wire [63:0] _GEN_69 = valid2_r & io_instRead_rvalid & ~reset_ic ? _GEN_63 : next_pc_r; // @[fetch.scala 233:64 fetch.scala 208:34]
  wire  _GEN_70 = valid2_r & io_instRead_rvalid & ~reset_ic ? _GEN_64 : wait_jmp_pc; // @[fetch.scala 233:64 fetch.scala 209:34]
  wire  _GEN_73 = excep2_r_en & valid2_r ? excep2_r_en : excep_buf_en; // @[fetch.scala 229:44 fetch.scala 230:23 fetch.scala 213:34]
  wire [127:0] _GEN_78 = excep2_r_en & valid2_r ? inst_buf : _GEN_66; // @[fetch.scala 229:44 fetch.scala 225:19]
  wire [1:0] _GEN_79 = excep2_r_en & valid2_r ? buf_bitmap : _GEN_67; // @[fetch.scala 229:44 fetch.scala 226:21]
  wire [63:0] _GEN_80 = excep2_r_en & valid2_r ? buf_start_pc : _GEN_68; // @[fetch.scala 229:44 fetch.scala 211:34]
  wire [63:0] _GEN_81 = excep2_r_en & valid2_r ? next_pc_r : _GEN_69; // @[fetch.scala 229:44 fetch.scala 208:34]
  wire  _GEN_82 = excep2_r_en & valid2_r ? wait_jmp_pc : _GEN_70; // @[fetch.scala 229:44 fetch.scala 209:34]
  wire  _GEN_85 = buf_bitmap == 2'h3 | excep_buf_en ? excep_buf_en : _GEN_73; // @[fetch.scala 228:49 fetch.scala 213:34]
  wire [127:0] _GEN_90 = buf_bitmap == 2'h3 | excep_buf_en ? inst_buf : _GEN_78; // @[fetch.scala 228:49 fetch.scala 225:19]
  wire [1:0] _GEN_91 = buf_bitmap == 2'h3 | excep_buf_en ? buf_bitmap : _GEN_79; // @[fetch.scala 228:49 fetch.scala 226:21]
  wire [63:0] _GEN_92 = buf_bitmap == 2'h3 | excep_buf_en ? buf_start_pc : _GEN_80; // @[fetch.scala 228:49 fetch.scala 211:34]
  wire [63:0] _GEN_93 = buf_bitmap == 2'h3 | excep_buf_en ? next_pc_r : _GEN_81; // @[fetch.scala 228:49 fetch.scala 208:34]
  wire  _GEN_94 = buf_bitmap == 2'h3 | excep_buf_en ? wait_jmp_pc : _GEN_82; // @[fetch.scala 228:49 fetch.scala 209:34]
  wire  _GEN_97 = _stall2_in_T & _GEN_85; // @[fetch.scala 227:20 fetch.scala 252:22]
  wire [127:0] next_inst_buf = _stall2_in_T ? _GEN_90 : inst_buf; // @[fetch.scala 227:20 fetch.scala 225:19]
  wire [1:0] next_buf_bitmap = _stall2_in_T ? _GEN_91 : buf_bitmap; // @[fetch.scala 227:20 fetch.scala 226:21]
  wire [63:0] _GEN_104 = _stall2_in_T ? _GEN_92 : buf_start_pc; // @[fetch.scala 227:20 fetch.scala 211:34]
  wire [63:0] _GEN_105 = _stall2_in_T ? _GEN_93 : next_pc_r; // @[fetch.scala 227:20 fetch.scala 208:34]
  wire  _GEN_106 = _stall2_in_T ? _GEN_94 : 1'h1; // @[fetch.scala 227:20 fetch.scala 254:21]
  wire [1:0] _GEN_107 = _stall2_in_T ? next_buf_bitmap : 2'h0; // @[fetch.scala 227:20 fetch.scala 248:20 fetch.scala 251:20]
  wire [127:0] _GEN_108 = _stall2_in_T ? next_inst_buf : inst_buf; // @[fetch.scala 227:20 fetch.scala 249:18 fetch.scala 210:34]
  wire [2:0] top_inst32_hi = buf_offset[2:0]; // @[fetch.scala 258:48]
  wire [5:0] _top_inst32_T = {top_inst32_hi,3'h0}; // @[Cat.scala 30:58]
  wire [127:0] top_inst32 = inst_buf >> _top_inst32_T; // @[fetch.scala 258:31]
  wire  _top_inst_T_1 = top_inst32[1:0] == 2'h3; // @[fetch.scala 262:41]
  wire [15:0] top_inst_lo = top_inst32[15:0]; // @[fetch.scala 262:87]
  wire [31:0] _top_inst_T_2 = {16'h0,top_inst_lo}; // @[Cat.scala 30:58]
  wire [127:0] _top_inst_T_3 = top_inst32[1:0] == 2'h3 ? top_inst32 : {{96'd0}, _top_inst_T_2}; // @[fetch.scala 262:24]
  wire  _T_22 = buf_bitmap == 2'h1; // @[fetch.scala 263:27]
  wire  _T_23 = buf_offset == 64'h6; // @[fetch.scala 264:25]
  wire  _T_27 = buf_offset <= 64'h4; // @[fetch.scala 267:31]
  wire [127:0] _GEN_111 = buf_offset <= 64'h4 ? _top_inst_T_3 : 128'h0; // @[fetch.scala 267:38 fetch.scala 269:22 fetch.scala 259:37]
  wire  _GEN_112 = buf_offset == 64'h6 & top_inst32[1:0] != 2'h3 | _T_27; // @[fetch.scala 264:60 fetch.scala 265:24]
  wire [127:0] _GEN_113 = buf_offset == 64'h6 & top_inst32[1:0] != 2'h3 ? {{96'd0}, _top_inst_T_2} : _GEN_111; // @[fetch.scala 264:60 fetch.scala 266:22]
  wire  _GEN_114 = buf_bitmap == 2'h1 & _GEN_112; // @[fetch.scala 263:35 fetch.scala 259:16]
  wire [127:0] _GEN_115 = buf_bitmap == 2'h1 ? _GEN_113 : 128'h0; // @[fetch.scala 263:35 fetch.scala 259:37]
  wire  inst_valid = _T_14 | _GEN_114; // @[fetch.scala 260:29 fetch.scala 261:20]
  wire [127:0] _GEN_117 = _T_14 ? _top_inst_T_3 : _GEN_115; // @[fetch.scala 260:29 fetch.scala 262:18]
  wire  fetch_page_fault_excep = excep_buf_cause == 64'hc; // @[fetch.scala 272:50]
  wire  cross_page_excep = fetch_page_fault_excep & _T_22 & _T_23 & _top_inst_T_1; // @[fetch.scala 273:95]
  wire [63:0] _excep3_r_T_tval = inst_valid ? 64'h0 : excep_buf_tval; // @[fetch.scala 277:31]
  wire [63:0] _excep3_r_T_pc = inst_valid ? 64'h0 : excep_buf_pc; // @[fetch.scala 277:31]
  wire [31:0] top_inst = _GEN_117[31:0]; // @[fetch.scala 257:24]
  wire [63:0] _excep3_r_tval_T_1 = next_pc_r + 64'h2; // @[fetch.scala 282:59]
  wire [63:0] _excep3_r_tval_T_2 = fetch_page_fault_excep ? next_pc_r : excep_buf_tval; // @[Mux.scala 47:69]
  wire [63:0] _excep3_r_tval_T_3 = cross_page_excep ? _excep3_r_tval_T_1 : _excep3_r_tval_T_2; // @[Mux.scala 47:69]
  wire [2:0] _next_pc_w_T_2 = top_inst[1:0] == 2'h3 ? 3'h4 : 3'h2; // @[fetch.scala 288:44]
  wire [63:0] _GEN_156 = {{61'd0}, _next_pc_w_T_2}; // @[fetch.scala 288:39]
  wire [63:0] next_pc_w = next_pc_r + _GEN_156; // @[fetch.scala 288:39]
  wire [63:0] _T_34 = next_pc_w - buf_start_pc; // @[fetch.scala 290:29]
  wire [63:0] _buf_start_pc_T_2 = buf_start_pc + 64'h8; // @[fetch.scala 291:46]
  wire [63:0] inst_buf_lo = next_inst_buf[127:64]; // @[fetch.scala 292:57]
  wire [127:0] _inst_buf_T = {64'h0,inst_buf_lo}; // @[Cat.scala 30:58]
  wire  buf_bitmap_lo = next_buf_bitmap[1]; // @[fetch.scala 293:60]
  wire [1:0] _buf_bitmap_T = {1'h0,buf_bitmap_lo}; // @[Cat.scala 30:58]
  wire  _T_38 = ~inst_valid; // @[fetch.scala 295:18]
  wire  _GEN_125 = hs_out ? 1'h0 : valid3_r; // @[fetch.scala 301:27 fetch.scala 302:22 fetch.scala 206:34]
  wire  _GEN_126 = (inst_valid | excep_buf_en) & (~valid3_r | hs_out) | _GEN_125; // @[fetch.scala 275:68 fetch.scala 276:25]
  wire  _GEN_139 = (inst_valid | excep_buf_en) & (~valid3_r | hs_out) & _T_38; // @[fetch.scala 275:68 fetch.scala 72:53]
  wire  _GEN_141 = _stall3_in_T & _GEN_126; // @[fetch.scala 274:25 fetch.scala 305:18]
  wire  _GEN_154 = _stall3_in_T & _GEN_139; // @[fetch.scala 274:25 fetch.scala 72:53]
  assign io_instRead_addr = hs1 ? io_va2pa_paddr : paddr2_r; // @[fetch.scala 201:28]
  assign io_instRead_arvalid = (hs1 | valid2_r) & _stall3_in_T & ~cur_excep_en; // @[fetch.scala 203:64]
  assign io_va2pa_vaddr = hs1 ? _cur_pc_T_1 : pc; // @[Mux.scala 47:69]
  assign io_va2pa_vvalid = hs_in & ~io_intr_in_en; // @[fetch.scala 150:30]
  assign io_if2id_inst = inst_r; // @[fetch.scala 308:25]
  assign io_if2id_pc = pc3_r; // @[fetch.scala 309:25]
  assign io_if2id_excep_cause = excep3_r_cause; // @[fetch.scala 310:25]
  assign io_if2id_excep_tval = excep3_r_tval; // @[fetch.scala 310:25]
  assign io_if2id_excep_en = excep3_r_en; // @[fetch.scala 310:25]
  assign io_if2id_excep_pc = excep3_r_pc; // @[fetch.scala 310:25]
  assign io_if2id_recov = recov3_r; // @[fetch.scala 312:25]
  assign io_if2id_valid = valid3_r; // @[fetch.scala 311:25]
  always @(posedge clock) begin
    if (reset) begin // @[fetch.scala 61:21]
      pc <= 64'h30000000; // @[fetch.scala 61:21]
    end else if (io_reg2if_valid) begin // @[Mux.scala 47:69]
      pc <= io_reg2if_seq_pc;
    end else if (io_wb2if_valid) begin // @[Mux.scala 47:69]
      pc <= io_wb2if_seq_pc;
    end else if (io_intr_in_en) begin // @[Mux.scala 47:69]
      pc <= cur_pc;
    end else begin
      pc <= _next_pc_T;
    end
    if (reset) begin // @[fetch.scala 63:26]
      drop1_r <= 1'h0; // @[fetch.scala 63:26]
    end else begin
      drop1_r <= _GEN_10;
    end
    if (reset) begin // @[fetch.scala 64:26]
      drop2_r <= 1'h0; // @[fetch.scala 64:26]
    end else begin
      drop2_r <= _GEN_54;
    end
    if (reset) begin // @[fetch.scala 65:26]
      drop3_r <= 1'h0; // @[fetch.scala 65:26]
    end else begin
      drop3_r <= _GEN_154;
    end
    if (reset) begin // @[fetch.scala 66:27]
      stall1_r <= 1'h0; // @[fetch.scala 66:27]
    end else begin
      stall1_r <= _GEN_10;
    end
    if (reset) begin // @[fetch.scala 67:27]
      stall2_r <= 1'h0; // @[fetch.scala 67:27]
    end else begin
      stall2_r <= _GEN_54;
    end
    if (reset) begin // @[fetch.scala 68:27]
      stall3_r <= 1'h0; // @[fetch.scala 68:27]
    end else begin
      stall3_r <= _GEN_154;
    end
    if (reset) begin // @[fetch.scala 71:27]
      recov3_r <= 1'h0; // @[fetch.scala 71:27]
    end else if (_stall3_in_T) begin // @[fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[fetch.scala 275:68]
        recov3_r <= _T_38;
      end
    end
    if (reset) begin // @[fetch.scala 91:24]
      state <= 1'h0; // @[fetch.scala 91:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      state <= _GEN_0;
    end else if (state) begin // @[Conditional.scala 39:67]
      if (drop1_in & ~stall1_in | io_recov) begin // @[fetch.scala 99:55]
        state <= 1'h0; // @[fetch.scala 100:23]
      end
    end
    if (reset) begin // @[fetch.scala 105:24]
      pc1_r <= 64'h0; // @[fetch.scala 105:24]
    end else if (hs1) begin // @[Mux.scala 47:69]
      pc1_r <= _cur_pc_T_1;
    end else begin
      pc1_r <= pc;
    end
    if (reset) begin // @[fetch.scala 107:30]
      excep1_r_cause <= 64'h0; // @[fetch.scala 107:30]
    end else if (hs_in) begin // @[fetch.scala 126:16]
      excep1_r_cause <= io_intr_in_cause; // @[fetch.scala 129:25]
    end
    if (reset) begin // @[fetch.scala 107:30]
      excep1_r_en <= 1'h0; // @[fetch.scala 107:30]
    end else if (hs_in) begin // @[fetch.scala 126:16]
      excep1_r_en <= io_intr_in_en; // @[fetch.scala 127:25]
    end
    if (reset) begin // @[fetch.scala 108:30]
      valid1_r <= 1'h0; // @[fetch.scala 108:30]
    end else begin
      valid1_r <= _GEN_14;
    end
    if (reset) begin // @[fetch.scala 156:30]
      valid2_r <= 1'h0; // @[fetch.scala 156:30]
    end else begin
      valid2_r <= _GEN_46;
    end
    if (reset) begin // @[fetch.scala 212:34]
      buf_bitmap <= 2'h0; // @[fetch.scala 212:34]
    end else if (_stall3_in_T) begin // @[fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[fetch.scala 275:68]
        if (_T_34 >= 64'h8 & buf_bitmap != 2'h0) begin // @[fetch.scala 290:74]
          buf_bitmap <= _buf_bitmap_T; // @[fetch.scala 293:28]
        end else begin
          buf_bitmap <= _GEN_107;
        end
      end else begin
        buf_bitmap <= _GEN_107;
      end
    end else begin
      buf_bitmap <= _GEN_107;
    end
    if (reset) begin // @[fetch.scala 213:34]
      excep_buf_en <= 1'h0; // @[fetch.scala 213:34]
    end else if (_stall3_in_T) begin // @[fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[fetch.scala 275:68]
        if (~inst_valid) begin // @[fetch.scala 295:30]
          excep_buf_en <= 1'h0; // @[fetch.scala 296:30]
        end else begin
          excep_buf_en <= _GEN_97;
        end
      end else begin
        excep_buf_en <= _GEN_97;
      end
    end else begin
      excep_buf_en <= _GEN_97;
    end
    if (reset) begin // @[fetch.scala 157:30]
      excep2_r_en <= 1'h0; // @[fetch.scala 157:30]
    end else if (_stall2_in_T) begin // @[fetch.scala 176:20]
      if (!(~hs1)) begin // @[fetch.scala 184:19]
        if (io_va2pa_pvalid) begin // @[fetch.scala 185:36]
          excep2_r_en <= 1'h0; // @[fetch.scala 187:28]
        end else begin
          excep2_r_en <= _GEN_24;
        end
      end
    end
    if (reset) begin // @[fetch.scala 217:30]
      reset_ic <= 1'h0; // @[fetch.scala 217:30]
    end else if (_stall2_in_T) begin // @[fetch.scala 227:20]
      if (io_instRead_rvalid) begin // @[fetch.scala 219:29]
        reset_ic <= 1'h0; // @[fetch.scala 220:18]
      end
    end else begin
      reset_ic <= reset_ic | valid2_r & ~excep2_r_en & ~io_instRead_rvalid; // @[fetch.scala 253:18]
    end
    if (reset) begin // @[fetch.scala 161:30]
      reset_tlb <= 1'h0; // @[fetch.scala 161:30]
    end else if (_stall2_in_T) begin // @[fetch.scala 176:20]
      if (_tlb_inp_valid_T_1) begin // @[fetch.scala 162:51]
        reset_tlb <= 1'h0; // @[fetch.scala 163:21]
      end
    end else begin
      reset_tlb <= ~_tlb_inp_valid_T_1; // @[fetch.scala 199:19]
    end
    if (reset) begin // @[fetch.scala 154:30]
      pc2_r <= 64'h0; // @[fetch.scala 154:30]
    end else if (_stall2_in_T) begin // @[fetch.scala 176:20]
      if (hs1) begin // @[fetch.scala 177:18]
        pc2_r <= pc1_r; // @[fetch.scala 179:29]
      end
    end
    if (reset) begin // @[fetch.scala 155:30]
      paddr2_r <= 32'h0; // @[fetch.scala 155:30]
    end else if (_stall2_in_T) begin // @[fetch.scala 176:20]
      if (!(~hs1)) begin // @[fetch.scala 184:19]
        if (io_va2pa_pvalid) begin // @[fetch.scala 185:36]
          paddr2_r <= io_va2pa_paddr; // @[fetch.scala 186:25]
        end
      end
    end
    if (reset) begin // @[fetch.scala 157:30]
      excep2_r_cause <= 64'h0; // @[fetch.scala 157:30]
    end else if (_stall2_in_T) begin // @[fetch.scala 176:20]
      if (!(~hs1)) begin // @[fetch.scala 184:19]
        if (!(io_va2pa_pvalid)) begin // @[fetch.scala 185:36]
          excep2_r_cause <= _GEN_26;
        end
      end
    end
    if (reset) begin // @[fetch.scala 157:30]
      excep2_r_tval <= 64'h0; // @[fetch.scala 157:30]
    end else if (_stall2_in_T) begin // @[fetch.scala 176:20]
      if (!(~hs1)) begin // @[fetch.scala 184:19]
        if (!(io_va2pa_pvalid)) begin // @[fetch.scala 185:36]
          excep2_r_tval <= _GEN_25;
        end
      end
    end
    if (reset) begin // @[fetch.scala 157:30]
      excep2_r_pc <= 64'h0; // @[fetch.scala 157:30]
    end else if (_stall2_in_T) begin // @[fetch.scala 176:20]
      if (!(~hs1)) begin // @[fetch.scala 184:19]
        if (!(io_va2pa_pvalid)) begin // @[fetch.scala 185:36]
          excep2_r_pc <= _GEN_23;
        end
      end
    end
    if (reset) begin // @[fetch.scala 205:34]
      pc3_r <= 64'h0; // @[fetch.scala 205:34]
    end else if (_stall3_in_T) begin // @[fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[fetch.scala 275:68]
        pc3_r <= next_pc_r; // @[fetch.scala 287:25]
      end
    end
    if (reset) begin // @[fetch.scala 206:34]
      valid3_r <= 1'h0; // @[fetch.scala 206:34]
    end else begin
      valid3_r <= _GEN_141;
    end
    if (reset) begin // @[fetch.scala 207:34]
      excep3_r_cause <= 64'h0; // @[fetch.scala 207:34]
    end else if (_stall3_in_T) begin // @[fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[fetch.scala 275:68]
        if (inst_valid) begin // @[fetch.scala 277:31]
          excep3_r_cause <= 64'h0;
        end else begin
          excep3_r_cause <= excep_buf_cause;
        end
      end
    end
    if (reset) begin // @[fetch.scala 207:34]
      excep3_r_tval <= 64'h0; // @[fetch.scala 207:34]
    end else if (_stall3_in_T) begin // @[fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[fetch.scala 275:68]
        if (update_excep_pc) begin // @[fetch.scala 279:34]
          excep3_r_tval <= _excep3_r_tval_T_3; // @[fetch.scala 281:31]
        end else begin
          excep3_r_tval <= _excep3_r_T_tval; // @[fetch.scala 277:25]
        end
      end
    end
    if (reset) begin // @[fetch.scala 207:34]
      excep3_r_en <= 1'h0; // @[fetch.scala 207:34]
    end else if (_stall3_in_T) begin // @[fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[fetch.scala 275:68]
        if (inst_valid) begin // @[fetch.scala 277:31]
          excep3_r_en <= 1'h0;
        end else begin
          excep3_r_en <= excep_buf_en;
        end
      end
    end
    if (reset) begin // @[fetch.scala 207:34]
      excep3_r_pc <= 64'h0; // @[fetch.scala 207:34]
    end else if (_stall3_in_T) begin // @[fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[fetch.scala 275:68]
        if (update_excep_pc) begin // @[fetch.scala 279:34]
          excep3_r_pc <= next_pc_r; // @[fetch.scala 280:29]
        end else begin
          excep3_r_pc <= _excep3_r_T_pc; // @[fetch.scala 277:25]
        end
      end
    end
    if (reset) begin // @[fetch.scala 208:34]
      next_pc_r <= 64'h0; // @[fetch.scala 208:34]
    end else if (_stall3_in_T) begin // @[fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[fetch.scala 275:68]
        next_pc_r <= next_pc_w; // @[fetch.scala 289:25]
      end else begin
        next_pc_r <= _GEN_105;
      end
    end else begin
      next_pc_r <= _GEN_105;
    end
    wait_jmp_pc <= reset | _GEN_106; // @[fetch.scala 209:34 fetch.scala 209:34]
    if (reset) begin // @[fetch.scala 210:34]
      inst_buf <= 128'h0; // @[fetch.scala 210:34]
    end else if (_stall3_in_T) begin // @[fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[fetch.scala 275:68]
        if (_T_34 >= 64'h8 & buf_bitmap != 2'h0) begin // @[fetch.scala 290:74]
          inst_buf <= _inst_buf_T; // @[fetch.scala 292:26]
        end else begin
          inst_buf <= _GEN_108;
        end
      end else begin
        inst_buf <= _GEN_108;
      end
    end else begin
      inst_buf <= _GEN_108;
    end
    if (reset) begin // @[fetch.scala 211:34]
      buf_start_pc <= 64'h0; // @[fetch.scala 211:34]
    end else if (_stall3_in_T) begin // @[fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[fetch.scala 275:68]
        if (_T_34 >= 64'h8 & buf_bitmap != 2'h0) begin // @[fetch.scala 290:74]
          buf_start_pc <= _buf_start_pc_T_2; // @[fetch.scala 291:30]
        end else begin
          buf_start_pc <= _GEN_104;
        end
      end else begin
        buf_start_pc <= _GEN_104;
      end
    end else begin
      buf_start_pc <= _GEN_104;
    end
    if (reset) begin // @[fetch.scala 213:34]
      excep_buf_cause <= 64'h0; // @[fetch.scala 213:34]
    end else if (_stall2_in_T) begin // @[fetch.scala 227:20]
      if (!(buf_bitmap == 2'h3 | excep_buf_en)) begin // @[fetch.scala 228:49]
        if (excep2_r_en & valid2_r) begin // @[fetch.scala 229:44]
          excep_buf_cause <= excep2_r_cause; // @[fetch.scala 230:23]
        end
      end
    end
    if (reset) begin // @[fetch.scala 213:34]
      excep_buf_tval <= 64'h0; // @[fetch.scala 213:34]
    end else if (_stall2_in_T) begin // @[fetch.scala 227:20]
      if (!(buf_bitmap == 2'h3 | excep_buf_en)) begin // @[fetch.scala 228:49]
        if (excep2_r_en & valid2_r) begin // @[fetch.scala 229:44]
          excep_buf_tval <= excep2_r_tval; // @[fetch.scala 230:23]
        end
      end
    end
    if (reset) begin // @[fetch.scala 213:34]
      excep_buf_pc <= 64'h0; // @[fetch.scala 213:34]
    end else if (_stall2_in_T) begin // @[fetch.scala 227:20]
      if (!(buf_bitmap == 2'h3 | excep_buf_en)) begin // @[fetch.scala 228:49]
        if (excep2_r_en & valid2_r) begin // @[fetch.scala 229:44]
          excep_buf_pc <= excep2_r_pc; // @[fetch.scala 230:23]
        end
      end
    end
    if (reset) begin // @[fetch.scala 214:34]
      inst_r <= 32'h0; // @[fetch.scala 214:34]
    end else if (_stall3_in_T) begin // @[fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[fetch.scala 275:68]
        if (inst_valid) begin // @[fetch.scala 278:31]
          inst_r <= top_inst;
        end else begin
          inst_r <= 32'h0;
        end
      end
    end
    if (reset) begin // @[fetch.scala 218:34]
      update_excep_pc <= 1'h0; // @[fetch.scala 218:34]
    end else if (_stall2_in_T) begin // @[fetch.scala 227:20]
      if (!(buf_bitmap == 2'h3 | excep_buf_en)) begin // @[fetch.scala 228:49]
        if (excep2_r_en & valid2_r) begin // @[fetch.scala 229:44]
          update_excep_pc <= ~wait_jmp_pc; // @[fetch.scala 232:29]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  drop1_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  drop2_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  drop3_r = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  stall1_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  stall2_r = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  stall3_r = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  recov3_r = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  pc1_r = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  excep1_r_cause = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  excep1_r_en = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  valid1_r = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  valid2_r = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  buf_bitmap = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  excep_buf_en = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  excep2_r_en = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  reset_ic = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  reset_tlb = _RAND_18[0:0];
  _RAND_19 = {2{`RANDOM}};
  pc2_r = _RAND_19[63:0];
  _RAND_20 = {1{`RANDOM}};
  paddr2_r = _RAND_20[31:0];
  _RAND_21 = {2{`RANDOM}};
  excep2_r_cause = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  excep2_r_tval = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  excep2_r_pc = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  pc3_r = _RAND_24[63:0];
  _RAND_25 = {1{`RANDOM}};
  valid3_r = _RAND_25[0:0];
  _RAND_26 = {2{`RANDOM}};
  excep3_r_cause = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  excep3_r_tval = _RAND_27[63:0];
  _RAND_28 = {1{`RANDOM}};
  excep3_r_en = _RAND_28[0:0];
  _RAND_29 = {2{`RANDOM}};
  excep3_r_pc = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  next_pc_r = _RAND_30[63:0];
  _RAND_31 = {1{`RANDOM}};
  wait_jmp_pc = _RAND_31[0:0];
  _RAND_32 = {4{`RANDOM}};
  inst_buf = _RAND_32[127:0];
  _RAND_33 = {2{`RANDOM}};
  buf_start_pc = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  excep_buf_cause = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  excep_buf_tval = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  excep_buf_pc = _RAND_36[63:0];
  _RAND_37 = {1{`RANDOM}};
  inst_r = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  update_excep_pc = _RAND_38[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_Decode(
  input         clock,
  input         reset,
  input  [31:0] io_if2id_inst,
  input  [63:0] io_if2id_pc,
  input  [63:0] io_if2id_excep_cause,
  input  [63:0] io_if2id_excep_tval,
  input         io_if2id_excep_en,
  input  [63:0] io_if2id_excep_pc,
  output        io_if2id_drop,
  output        io_if2id_stall,
  input         io_if2id_recov,
  input         io_if2id_valid,
  output        io_if2id_ready,
  output [31:0] io_id2df_inst,
  output [63:0] io_id2df_pc,
  output [63:0] io_id2df_excep_cause,
  output [63:0] io_id2df_excep_tval,
  output        io_id2df_excep_en,
  output [63:0] io_id2df_excep_pc,
  output [1:0]  io_id2df_excep_etype,
  output [4:0]  io_id2df_ctrl_aluOp,
  output        io_id2df_ctrl_aluWidth,
  output [4:0]  io_id2df_ctrl_dcMode,
  output        io_id2df_ctrl_writeRegEn,
  output        io_id2df_ctrl_writeCSREn,
  output [2:0]  io_id2df_ctrl_brType,
  output [4:0]  io_id2df_rs1,
  output        io_id2df_rrs1,
  output [63:0] io_id2df_rs1_d,
  output [11:0] io_id2df_rs2,
  output        io_id2df_rrs2,
  output [63:0] io_id2df_rs2_d,
  output [4:0]  io_id2df_dst,
  output [63:0] io_id2df_dst_d,
  output [1:0]  io_id2df_jmp_type,
  output [1:0]  io_id2df_special,
  output [5:0]  io_id2df_swap,
  output [1:0]  io_id2df_indi,
  input         io_id2df_drop,
  input         io_id2df_stall,
  output        io_id2df_recov,
  output        io_id2df_valid,
  input         io_id2df_ready,
  input  [1:0]  io_idState_priv
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  reg  drop_r; // @[decode.scala 17:30]
  reg  stall_r; // @[decode.scala 18:30]
  wire  drop_in = drop_r | io_id2df_drop; // @[decode.scala 20:30]
  wire  _io_if2id_stall_T = ~io_id2df_drop; // @[decode.scala 22:36]
  reg [31:0] inst_r; // @[decode.scala 23:30]
  reg [63:0] pc_r; // @[decode.scala 24:30]
  reg [63:0] excep_r_cause; // @[decode.scala 25:30]
  reg [63:0] excep_r_tval; // @[decode.scala 25:30]
  reg  excep_r_en; // @[decode.scala 25:30]
  reg [63:0] excep_r_pc; // @[decode.scala 25:30]
  reg [1:0] excep_r_etype; // @[decode.scala 25:30]
  reg [4:0] ctrl_r_aluOp; // @[decode.scala 26:30]
  reg  ctrl_r_aluWidth; // @[decode.scala 26:30]
  reg [4:0] ctrl_r_dcMode; // @[decode.scala 26:30]
  reg  ctrl_r_writeRegEn; // @[decode.scala 26:30]
  reg  ctrl_r_writeCSREn; // @[decode.scala 26:30]
  reg [2:0] ctrl_r_brType; // @[decode.scala 26:30]
  reg [4:0] rs1_r; // @[decode.scala 27:30]
  reg  rrs1_r; // @[decode.scala 28:30]
  reg [63:0] rs1_d_r; // @[decode.scala 29:30]
  reg [11:0] rs2_r; // @[decode.scala 30:30]
  reg  rrs2_r; // @[decode.scala 31:30]
  reg [63:0] rs2_d_r; // @[decode.scala 32:30]
  reg [4:0] dst_r; // @[decode.scala 33:30]
  reg [63:0] dst_d_r; // @[decode.scala 34:30]
  reg [1:0] jmp_type_r; // @[decode.scala 35:30]
  reg [1:0] special_r; // @[decode.scala 36:30]
  reg [5:0] swap_r; // @[decode.scala 37:30]
  reg [1:0] indi_r; // @[decode.scala 38:30]
  reg  recov_r; // @[decode.scala 39:30]
  reg  valid_r; // @[decode.scala 40:30]
  wire  hs_out = io_id2df_ready & io_id2df_valid; // @[decode.scala 46:33]
  wire  hs_in = io_if2id_ready & io_if2id_valid; // @[decode.scala 47:33]
  wire [31:0] _instType_T = io_if2id_inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _instType_T_1 = 32'h37 == _instType_T; // @[Lookup.scala 31:38]
  wire  _instType_T_3 = 32'h17 == _instType_T; // @[Lookup.scala 31:38]
  wire  _instType_T_5 = 32'h6f == _instType_T; // @[Lookup.scala 31:38]
  wire [31:0] _instType_T_6 = io_if2id_inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _instType_T_7 = 32'h67 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_9 = 32'h63 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_11 = 32'h1063 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_13 = 32'h4063 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_15 = 32'h5063 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_17 = 32'h6063 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_19 = 32'h7063 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_21 = 32'h3 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_23 = 32'h1003 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_25 = 32'h2003 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_27 = 32'h3003 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_29 = 32'h4003 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_31 = 32'h5003 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_33 = 32'h6003 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_35 = 32'h23 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_37 = 32'h1023 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_39 = 32'h2023 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_41 = 32'h3023 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_43 = 32'h13 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_45 = 32'h2013 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_47 = 32'h3013 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_49 = 32'h4013 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_51 = 32'h6013 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_53 = 32'h7013 == _instType_T_6; // @[Lookup.scala 31:38]
  wire [31:0] _instType_T_54 = io_if2id_inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _instType_T_55 = 32'h1013 == _instType_T_54; // @[Lookup.scala 31:38]
  wire  _instType_T_57 = 32'h5013 == _instType_T_54; // @[Lookup.scala 31:38]
  wire  _instType_T_59 = 32'h40005013 == _instType_T_54; // @[Lookup.scala 31:38]
  wire [31:0] _instType_T_60 = io_if2id_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _instType_T_61 = 32'h33 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_63 = 32'h40000033 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_65 = 32'h1033 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_67 = 32'h2033 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_69 = 32'h3033 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_71 = 32'h4033 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_73 = 32'h5033 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_75 = 32'h40005033 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_77 = 32'h6033 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_79 = 32'h7033 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_81 = 32'h2000033 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_83 = 32'h2001033 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_85 = 32'h2003033 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_87 = 32'h2002033 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_89 = 32'h2004033 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_91 = 32'h2005033 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_93 = 32'h2006033 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_95 = 32'h2007033 == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_97 = 32'h200003b == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_99 = 32'h200403b == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_101 = 32'h200503b == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_103 = 32'h200603b == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_105 = 32'h200703b == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_107 = 32'h1b == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_109 = 32'h101b == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_111 = 32'h501b == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_113 = 32'h4000501b == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_115 = 32'h3b == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_117 = 32'h4000003b == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_119 = 32'h103b == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_121 = 32'h503b == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_123 = 32'h4000503b == _instType_T_60; // @[Lookup.scala 31:38]
  wire  _instType_T_125 = 32'h1073 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_127 = 32'h2073 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_129 = 32'h3073 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_131 = 32'h5073 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_133 = 32'h6073 == _instType_T_6; // @[Lookup.scala 31:38]
  wire  _instType_T_135 = 32'h7073 == _instType_T_6; // @[Lookup.scala 31:38]
  wire [31:0] _instType_T_136 = io_if2id_inst & 32'hf9f0707f; // @[Lookup.scala 31:38]
  wire  _instType_T_137 = 32'h1000202f == _instType_T_136; // @[Lookup.scala 31:38]
  wire [31:0] _instType_T_138 = io_if2id_inst & 32'hf800707f; // @[Lookup.scala 31:38]
  wire  _instType_T_139 = 32'h1800202f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_141 = 32'h800202f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_143 = 32'h202f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_145 = 32'h2000202f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_147 = 32'h6000202f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_149 = 32'h4000202f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_151 = 32'h8000202f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_153 = 32'ha000202f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_155 = 32'hc000202f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_157 = 32'he000202f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_159 = 32'h1000302f == _instType_T_136; // @[Lookup.scala 31:38]
  wire  _instType_T_161 = 32'h1800302f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_163 = 32'h800302f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_165 = 32'h302f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_167 = 32'h4000302f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_169 = 32'h2000302f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_171 = 32'h6000302f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_173 = 32'h8000302f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_175 = 32'ha000302f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_177 = 32'hc000302f == _instType_T_138; // @[Lookup.scala 31:38]
  wire  _instType_T_179 = 32'he000302f == _instType_T_138; // @[Lookup.scala 31:38]
  wire [31:0] _instType_T_180 = io_if2id_inst & 32'hf00fffff; // @[Lookup.scala 31:38]
  wire  _instType_T_181 = 32'hf == _instType_T_180; // @[Lookup.scala 31:38]
  wire  _instType_T_183 = 32'h100f == io_if2id_inst; // @[Lookup.scala 31:38]
  wire [31:0] _instType_T_184 = io_if2id_inst & 32'hfe007fff; // @[Lookup.scala 31:38]
  wire  _instType_T_185 = 32'h12000073 == _instType_T_184; // @[Lookup.scala 31:38]
  wire  _instType_T_187 = 32'h10500073 == io_if2id_inst; // @[Lookup.scala 31:38]
  wire  _instType_T_189 = 32'h6b == io_if2id_inst; // @[Lookup.scala 31:38]
  wire [2:0] _instType_T_190 = _instType_T_189 ? 3'h0 : 3'h7; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_191 = _instType_T_187 ? 3'h0 : _instType_T_190; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_192 = _instType_T_185 ? 3'h0 : _instType_T_191; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_193 = _instType_T_183 ? 3'h0 : _instType_T_192; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_194 = _instType_T_181 ? 3'h0 : _instType_T_193; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_195 = _instType_T_179 ? 3'h1 : _instType_T_194; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_196 = _instType_T_177 ? 3'h1 : _instType_T_195; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_197 = _instType_T_175 ? 3'h1 : _instType_T_196; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_198 = _instType_T_173 ? 3'h1 : _instType_T_197; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_199 = _instType_T_171 ? 3'h1 : _instType_T_198; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_200 = _instType_T_169 ? 3'h1 : _instType_T_199; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_201 = _instType_T_167 ? 3'h1 : _instType_T_200; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_202 = _instType_T_165 ? 3'h1 : _instType_T_201; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_203 = _instType_T_163 ? 3'h1 : _instType_T_202; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_204 = _instType_T_161 ? 3'h1 : _instType_T_203; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_205 = _instType_T_159 ? 3'h1 : _instType_T_204; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_206 = _instType_T_157 ? 3'h1 : _instType_T_205; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_207 = _instType_T_155 ? 3'h1 : _instType_T_206; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_208 = _instType_T_153 ? 3'h1 : _instType_T_207; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_209 = _instType_T_151 ? 3'h1 : _instType_T_208; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_210 = _instType_T_149 ? 3'h1 : _instType_T_209; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_211 = _instType_T_147 ? 3'h1 : _instType_T_210; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_212 = _instType_T_145 ? 3'h1 : _instType_T_211; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_213 = _instType_T_143 ? 3'h1 : _instType_T_212; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_214 = _instType_T_141 ? 3'h1 : _instType_T_213; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_215 = _instType_T_139 ? 3'h1 : _instType_T_214; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_216 = _instType_T_137 ? 3'h1 : _instType_T_215; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_217 = _instType_T_135 ? 3'h2 : _instType_T_216; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_218 = _instType_T_133 ? 3'h2 : _instType_T_217; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_219 = _instType_T_131 ? 3'h2 : _instType_T_218; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_220 = _instType_T_129 ? 3'h2 : _instType_T_219; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_221 = _instType_T_127 ? 3'h2 : _instType_T_220; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_222 = _instType_T_125 ? 3'h2 : _instType_T_221; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_223 = _instType_T_123 ? 3'h1 : _instType_T_222; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_224 = _instType_T_121 ? 3'h1 : _instType_T_223; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_225 = _instType_T_119 ? 3'h1 : _instType_T_224; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_226 = _instType_T_117 ? 3'h1 : _instType_T_225; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_227 = _instType_T_115 ? 3'h1 : _instType_T_226; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_228 = _instType_T_113 ? 3'h2 : _instType_T_227; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_229 = _instType_T_111 ? 3'h2 : _instType_T_228; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_230 = _instType_T_109 ? 3'h2 : _instType_T_229; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_231 = _instType_T_107 ? 3'h2 : _instType_T_230; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_232 = _instType_T_105 ? 3'h1 : _instType_T_231; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_233 = _instType_T_103 ? 3'h1 : _instType_T_232; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_234 = _instType_T_101 ? 3'h1 : _instType_T_233; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_235 = _instType_T_99 ? 3'h1 : _instType_T_234; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_236 = _instType_T_97 ? 3'h1 : _instType_T_235; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_237 = _instType_T_95 ? 3'h1 : _instType_T_236; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_238 = _instType_T_93 ? 3'h1 : _instType_T_237; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_239 = _instType_T_91 ? 3'h1 : _instType_T_238; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_240 = _instType_T_89 ? 3'h1 : _instType_T_239; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_241 = _instType_T_87 ? 3'h1 : _instType_T_240; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_242 = _instType_T_85 ? 3'h1 : _instType_T_241; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_243 = _instType_T_83 ? 3'h1 : _instType_T_242; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_244 = _instType_T_81 ? 3'h1 : _instType_T_243; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_245 = _instType_T_79 ? 3'h1 : _instType_T_244; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_246 = _instType_T_77 ? 3'h1 : _instType_T_245; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_247 = _instType_T_75 ? 3'h1 : _instType_T_246; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_248 = _instType_T_73 ? 3'h1 : _instType_T_247; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_249 = _instType_T_71 ? 3'h1 : _instType_T_248; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_250 = _instType_T_69 ? 3'h1 : _instType_T_249; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_251 = _instType_T_67 ? 3'h1 : _instType_T_250; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_252 = _instType_T_65 ? 3'h1 : _instType_T_251; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_253 = _instType_T_63 ? 3'h1 : _instType_T_252; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_254 = _instType_T_61 ? 3'h1 : _instType_T_253; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_255 = _instType_T_59 ? 3'h2 : _instType_T_254; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_256 = _instType_T_57 ? 3'h2 : _instType_T_255; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_257 = _instType_T_55 ? 3'h2 : _instType_T_256; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_258 = _instType_T_53 ? 3'h2 : _instType_T_257; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_259 = _instType_T_51 ? 3'h2 : _instType_T_258; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_260 = _instType_T_49 ? 3'h2 : _instType_T_259; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_261 = _instType_T_47 ? 3'h2 : _instType_T_260; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_262 = _instType_T_45 ? 3'h2 : _instType_T_261; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_263 = _instType_T_43 ? 3'h2 : _instType_T_262; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_264 = _instType_T_41 ? 3'h3 : _instType_T_263; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_265 = _instType_T_39 ? 3'h3 : _instType_T_264; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_266 = _instType_T_37 ? 3'h3 : _instType_T_265; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_267 = _instType_T_35 ? 3'h3 : _instType_T_266; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_268 = _instType_T_33 ? 3'h2 : _instType_T_267; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_269 = _instType_T_31 ? 3'h2 : _instType_T_268; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_270 = _instType_T_29 ? 3'h2 : _instType_T_269; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_271 = _instType_T_27 ? 3'h2 : _instType_T_270; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_272 = _instType_T_25 ? 3'h2 : _instType_T_271; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_273 = _instType_T_23 ? 3'h2 : _instType_T_272; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_274 = _instType_T_21 ? 3'h2 : _instType_T_273; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_275 = _instType_T_19 ? 3'h4 : _instType_T_274; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_276 = _instType_T_17 ? 3'h4 : _instType_T_275; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_277 = _instType_T_15 ? 3'h4 : _instType_T_276; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_278 = _instType_T_13 ? 3'h4 : _instType_T_277; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_279 = _instType_T_11 ? 3'h4 : _instType_T_278; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_280 = _instType_T_9 ? 3'h4 : _instType_T_279; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_281 = _instType_T_7 ? 3'h2 : _instType_T_280; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_282 = _instType_T_5 ? 3'h6 : _instType_T_281; // @[Lookup.scala 33:37]
  wire [2:0] _instType_T_283 = _instType_T_3 ? 3'h5 : _instType_T_282; // @[Lookup.scala 33:37]
  wire [2:0] dType = _instType_T_1 ? 3'h5 : _instType_T_283; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_289 = _instType_T_179 ? 5'h1 : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_290 = _instType_T_177 ? 5'h1 : _instType_T_289; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_291 = _instType_T_175 ? 5'h1 : _instType_T_290; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_292 = _instType_T_173 ? 5'h1 : _instType_T_291; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_293 = _instType_T_171 ? 5'h1 : _instType_T_292; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_294 = _instType_T_169 ? 5'h1 : _instType_T_293; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_295 = _instType_T_167 ? 5'h1 : _instType_T_294; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_296 = _instType_T_165 ? 5'h1 : _instType_T_295; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_297 = _instType_T_163 ? 5'h1 : _instType_T_296; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_298 = _instType_T_161 ? 5'h1 : _instType_T_297; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_299 = _instType_T_159 ? 5'h1 : _instType_T_298; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_300 = _instType_T_157 ? 5'h1 : _instType_T_299; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_301 = _instType_T_155 ? 5'h1 : _instType_T_300; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_302 = _instType_T_153 ? 5'h1 : _instType_T_301; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_303 = _instType_T_151 ? 5'h1 : _instType_T_302; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_304 = _instType_T_149 ? 5'h1 : _instType_T_303; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_305 = _instType_T_147 ? 5'h1 : _instType_T_304; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_306 = _instType_T_145 ? 5'h1 : _instType_T_305; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_307 = _instType_T_143 ? 5'h1 : _instType_T_306; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_308 = _instType_T_141 ? 5'h1 : _instType_T_307; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_309 = _instType_T_139 ? 5'h1 : _instType_T_308; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_310 = _instType_T_137 ? 5'h1 : _instType_T_309; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_311 = _instType_T_135 ? 5'h15 : _instType_T_310; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_312 = _instType_T_133 ? 5'h5 : _instType_T_311; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_313 = _instType_T_131 ? 5'h1 : _instType_T_312; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_314 = _instType_T_129 ? 5'h15 : _instType_T_313; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_315 = _instType_T_127 ? 5'h5 : _instType_T_314; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_316 = _instType_T_125 ? 5'h1 : _instType_T_315; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_317 = _instType_T_123 ? 5'h9 : _instType_T_316; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_318 = _instType_T_121 ? 5'h8 : _instType_T_317; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_319 = _instType_T_119 ? 5'h7 : _instType_T_318; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_320 = _instType_T_117 ? 5'ha : _instType_T_319; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_321 = _instType_T_115 ? 5'h3 : _instType_T_320; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_322 = _instType_T_113 ? 5'h9 : _instType_T_321; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_323 = _instType_T_111 ? 5'h8 : _instType_T_322; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_324 = _instType_T_109 ? 5'h7 : _instType_T_323; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_325 = _instType_T_107 ? 5'h3 : _instType_T_324; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_326 = _instType_T_105 ? 5'h14 : _instType_T_325; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_327 = _instType_T_103 ? 5'h13 : _instType_T_326; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_328 = _instType_T_101 ? 5'h12 : _instType_T_327; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_329 = _instType_T_99 ? 5'h11 : _instType_T_328; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_330 = _instType_T_97 ? 5'hd : _instType_T_329; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_331 = _instType_T_95 ? 5'h14 : _instType_T_330; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_332 = _instType_T_93 ? 5'h13 : _instType_T_331; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_333 = _instType_T_91 ? 5'h12 : _instType_T_332; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_334 = _instType_T_89 ? 5'h11 : _instType_T_333; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_335 = _instType_T_87 ? 5'h10 : _instType_T_334; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_336 = _instType_T_85 ? 5'hf : _instType_T_335; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_337 = _instType_T_83 ? 5'he : _instType_T_336; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_338 = _instType_T_81 ? 5'hd : _instType_T_337; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_339 = _instType_T_79 ? 5'h6 : _instType_T_338; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_340 = _instType_T_77 ? 5'h5 : _instType_T_339; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_341 = _instType_T_75 ? 5'h9 : _instType_T_340; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_342 = _instType_T_73 ? 5'h8 : _instType_T_341; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_343 = _instType_T_71 ? 5'h4 : _instType_T_342; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_344 = _instType_T_69 ? 5'hc : _instType_T_343; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_345 = _instType_T_67 ? 5'hb : _instType_T_344; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_346 = _instType_T_65 ? 5'h7 : _instType_T_345; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_347 = _instType_T_63 ? 5'ha : _instType_T_346; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_348 = _instType_T_61 ? 5'h3 : _instType_T_347; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_349 = _instType_T_59 ? 5'h9 : _instType_T_348; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_350 = _instType_T_57 ? 5'h8 : _instType_T_349; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_351 = _instType_T_55 ? 5'h7 : _instType_T_350; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_352 = _instType_T_53 ? 5'h6 : _instType_T_351; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_353 = _instType_T_51 ? 5'h5 : _instType_T_352; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_354 = _instType_T_49 ? 5'h4 : _instType_T_353; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_355 = _instType_T_47 ? 5'hc : _instType_T_354; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_356 = _instType_T_45 ? 5'hb : _instType_T_355; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_357 = _instType_T_43 ? 5'h3 : _instType_T_356; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_358 = _instType_T_41 ? 5'h3 : _instType_T_357; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_359 = _instType_T_39 ? 5'h3 : _instType_T_358; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_360 = _instType_T_37 ? 5'h3 : _instType_T_359; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_361 = _instType_T_35 ? 5'h3 : _instType_T_360; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_362 = _instType_T_33 ? 5'h3 : _instType_T_361; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_363 = _instType_T_31 ? 5'h3 : _instType_T_362; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_364 = _instType_T_29 ? 5'h3 : _instType_T_363; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_365 = _instType_T_27 ? 5'h3 : _instType_T_364; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_366 = _instType_T_25 ? 5'h3 : _instType_T_365; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_367 = _instType_T_23 ? 5'h3 : _instType_T_366; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_368 = _instType_T_21 ? 5'h3 : _instType_T_367; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_369 = _instType_T_19 ? 5'h0 : _instType_T_368; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_370 = _instType_T_17 ? 5'h0 : _instType_T_369; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_371 = _instType_T_15 ? 5'h0 : _instType_T_370; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_372 = _instType_T_13 ? 5'h0 : _instType_T_371; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_373 = _instType_T_11 ? 5'h0 : _instType_T_372; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_374 = _instType_T_9 ? 5'h0 : _instType_T_373; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_375 = _instType_T_7 ? 5'h2 : _instType_T_374; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_376 = _instType_T_5 ? 5'h2 : _instType_T_375; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_377 = _instType_T_3 ? 5'h3 : _instType_T_376; // @[Lookup.scala 33:37]
  wire [4:0] instType_1 = _instType_T_1 ? 5'h1 : _instType_T_377; // @[Lookup.scala 33:37]
  wire  _instType_T_425 = _instType_T_95 ? 1'h0 : _instType_T_97 | (_instType_T_99 | (_instType_T_101 | (_instType_T_103
     | (_instType_T_105 | (_instType_T_107 | (_instType_T_109 | (_instType_T_111 | (_instType_T_113 | (_instType_T_115
     | (_instType_T_117 | (_instType_T_119 | (_instType_T_121 | _instType_T_123)))))))))))); // @[Lookup.scala 33:37]
  wire  _instType_T_426 = _instType_T_93 ? 1'h0 : _instType_T_425; // @[Lookup.scala 33:37]
  wire  _instType_T_427 = _instType_T_91 ? 1'h0 : _instType_T_426; // @[Lookup.scala 33:37]
  wire  _instType_T_428 = _instType_T_89 ? 1'h0 : _instType_T_427; // @[Lookup.scala 33:37]
  wire  _instType_T_429 = _instType_T_87 ? 1'h0 : _instType_T_428; // @[Lookup.scala 33:37]
  wire  _instType_T_430 = _instType_T_85 ? 1'h0 : _instType_T_429; // @[Lookup.scala 33:37]
  wire  _instType_T_431 = _instType_T_83 ? 1'h0 : _instType_T_430; // @[Lookup.scala 33:37]
  wire  _instType_T_432 = _instType_T_81 ? 1'h0 : _instType_T_431; // @[Lookup.scala 33:37]
  wire  _instType_T_433 = _instType_T_79 ? 1'h0 : _instType_T_432; // @[Lookup.scala 33:37]
  wire  _instType_T_434 = _instType_T_77 ? 1'h0 : _instType_T_433; // @[Lookup.scala 33:37]
  wire  _instType_T_435 = _instType_T_75 ? 1'h0 : _instType_T_434; // @[Lookup.scala 33:37]
  wire  _instType_T_436 = _instType_T_73 ? 1'h0 : _instType_T_435; // @[Lookup.scala 33:37]
  wire  _instType_T_437 = _instType_T_71 ? 1'h0 : _instType_T_436; // @[Lookup.scala 33:37]
  wire  _instType_T_438 = _instType_T_69 ? 1'h0 : _instType_T_437; // @[Lookup.scala 33:37]
  wire  _instType_T_439 = _instType_T_67 ? 1'h0 : _instType_T_438; // @[Lookup.scala 33:37]
  wire  _instType_T_440 = _instType_T_65 ? 1'h0 : _instType_T_439; // @[Lookup.scala 33:37]
  wire  _instType_T_441 = _instType_T_63 ? 1'h0 : _instType_T_440; // @[Lookup.scala 33:37]
  wire  _instType_T_442 = _instType_T_61 ? 1'h0 : _instType_T_441; // @[Lookup.scala 33:37]
  wire  _instType_T_443 = _instType_T_59 ? 1'h0 : _instType_T_442; // @[Lookup.scala 33:37]
  wire  _instType_T_444 = _instType_T_57 ? 1'h0 : _instType_T_443; // @[Lookup.scala 33:37]
  wire  _instType_T_445 = _instType_T_55 ? 1'h0 : _instType_T_444; // @[Lookup.scala 33:37]
  wire  _instType_T_446 = _instType_T_53 ? 1'h0 : _instType_T_445; // @[Lookup.scala 33:37]
  wire  _instType_T_447 = _instType_T_51 ? 1'h0 : _instType_T_446; // @[Lookup.scala 33:37]
  wire  _instType_T_448 = _instType_T_49 ? 1'h0 : _instType_T_447; // @[Lookup.scala 33:37]
  wire  _instType_T_449 = _instType_T_47 ? 1'h0 : _instType_T_448; // @[Lookup.scala 33:37]
  wire  _instType_T_450 = _instType_T_45 ? 1'h0 : _instType_T_449; // @[Lookup.scala 33:37]
  wire  _instType_T_451 = _instType_T_43 ? 1'h0 : _instType_T_450; // @[Lookup.scala 33:37]
  wire  _instType_T_452 = _instType_T_41 ? 1'h0 : _instType_T_451; // @[Lookup.scala 33:37]
  wire  _instType_T_453 = _instType_T_39 ? 1'h0 : _instType_T_452; // @[Lookup.scala 33:37]
  wire  _instType_T_454 = _instType_T_37 ? 1'h0 : _instType_T_453; // @[Lookup.scala 33:37]
  wire  _instType_T_455 = _instType_T_35 ? 1'h0 : _instType_T_454; // @[Lookup.scala 33:37]
  wire  _instType_T_456 = _instType_T_33 ? 1'h0 : _instType_T_455; // @[Lookup.scala 33:37]
  wire  _instType_T_457 = _instType_T_31 ? 1'h0 : _instType_T_456; // @[Lookup.scala 33:37]
  wire  _instType_T_458 = _instType_T_29 ? 1'h0 : _instType_T_457; // @[Lookup.scala 33:37]
  wire  _instType_T_459 = _instType_T_27 ? 1'h0 : _instType_T_458; // @[Lookup.scala 33:37]
  wire  _instType_T_460 = _instType_T_25 ? 1'h0 : _instType_T_459; // @[Lookup.scala 33:37]
  wire  _instType_T_461 = _instType_T_23 ? 1'h0 : _instType_T_460; // @[Lookup.scala 33:37]
  wire  _instType_T_462 = _instType_T_21 ? 1'h0 : _instType_T_461; // @[Lookup.scala 33:37]
  wire  _instType_T_463 = _instType_T_19 ? 1'h0 : _instType_T_462; // @[Lookup.scala 33:37]
  wire  _instType_T_464 = _instType_T_17 ? 1'h0 : _instType_T_463; // @[Lookup.scala 33:37]
  wire  _instType_T_465 = _instType_T_15 ? 1'h0 : _instType_T_464; // @[Lookup.scala 33:37]
  wire  _instType_T_466 = _instType_T_13 ? 1'h0 : _instType_T_465; // @[Lookup.scala 33:37]
  wire  _instType_T_467 = _instType_T_11 ? 1'h0 : _instType_T_466; // @[Lookup.scala 33:37]
  wire  _instType_T_468 = _instType_T_9 ? 1'h0 : _instType_T_467; // @[Lookup.scala 33:37]
  wire  _instType_T_469 = _instType_T_7 ? 1'h0 : _instType_T_468; // @[Lookup.scala 33:37]
  wire  _instType_T_470 = _instType_T_5 ? 1'h0 : _instType_T_469; // @[Lookup.scala 33:37]
  wire  _instType_T_471 = _instType_T_3 ? 1'h0 : _instType_T_470; // @[Lookup.scala 33:37]
  wire  instType_2 = _instType_T_1 ? 1'h0 : _instType_T_471; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_477 = _instType_T_179 ? 5'hf : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_478 = _instType_T_177 ? 5'hf : _instType_T_477; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_479 = _instType_T_175 ? 5'hf : _instType_T_478; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_480 = _instType_T_173 ? 5'hf : _instType_T_479; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_481 = _instType_T_171 ? 5'hf : _instType_T_480; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_482 = _instType_T_169 ? 5'hf : _instType_T_481; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_483 = _instType_T_167 ? 5'hf : _instType_T_482; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_484 = _instType_T_165 ? 5'hf : _instType_T_483; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_485 = _instType_T_163 ? 5'hf : _instType_T_484; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_486 = _instType_T_161 ? 5'hb : _instType_T_485; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_487 = _instType_T_159 ? 5'h7 : _instType_T_486; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_488 = _instType_T_157 ? 5'he : _instType_T_487; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_489 = _instType_T_155 ? 5'he : _instType_T_488; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_490 = _instType_T_153 ? 5'he : _instType_T_489; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_491 = _instType_T_151 ? 5'he : _instType_T_490; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_492 = _instType_T_149 ? 5'he : _instType_T_491; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_493 = _instType_T_147 ? 5'he : _instType_T_492; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_494 = _instType_T_145 ? 5'he : _instType_T_493; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_495 = _instType_T_143 ? 5'he : _instType_T_494; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_496 = _instType_T_141 ? 5'he : _instType_T_495; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_497 = _instType_T_139 ? 5'ha : _instType_T_496; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_498 = _instType_T_137 ? 5'h6 : _instType_T_497; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_499 = _instType_T_135 ? 5'h0 : _instType_T_498; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_500 = _instType_T_133 ? 5'h0 : _instType_T_499; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_501 = _instType_T_131 ? 5'h0 : _instType_T_500; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_502 = _instType_T_129 ? 5'h0 : _instType_T_501; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_503 = _instType_T_127 ? 5'h0 : _instType_T_502; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_504 = _instType_T_125 ? 5'h0 : _instType_T_503; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_505 = _instType_T_123 ? 5'h0 : _instType_T_504; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_506 = _instType_T_121 ? 5'h0 : _instType_T_505; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_507 = _instType_T_119 ? 5'h0 : _instType_T_506; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_508 = _instType_T_117 ? 5'h0 : _instType_T_507; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_509 = _instType_T_115 ? 5'h0 : _instType_T_508; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_510 = _instType_T_113 ? 5'h0 : _instType_T_509; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_511 = _instType_T_111 ? 5'h0 : _instType_T_510; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_512 = _instType_T_109 ? 5'h0 : _instType_T_511; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_513 = _instType_T_107 ? 5'h0 : _instType_T_512; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_514 = _instType_T_105 ? 5'h0 : _instType_T_513; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_515 = _instType_T_103 ? 5'h0 : _instType_T_514; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_516 = _instType_T_101 ? 5'h0 : _instType_T_515; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_517 = _instType_T_99 ? 5'h0 : _instType_T_516; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_518 = _instType_T_97 ? 5'h0 : _instType_T_517; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_519 = _instType_T_95 ? 5'h0 : _instType_T_518; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_520 = _instType_T_93 ? 5'h0 : _instType_T_519; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_521 = _instType_T_91 ? 5'h0 : _instType_T_520; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_522 = _instType_T_89 ? 5'h0 : _instType_T_521; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_523 = _instType_T_87 ? 5'h0 : _instType_T_522; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_524 = _instType_T_85 ? 5'h0 : _instType_T_523; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_525 = _instType_T_83 ? 5'h0 : _instType_T_524; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_526 = _instType_T_81 ? 5'h0 : _instType_T_525; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_527 = _instType_T_79 ? 5'h0 : _instType_T_526; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_528 = _instType_T_77 ? 5'h0 : _instType_T_527; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_529 = _instType_T_75 ? 5'h0 : _instType_T_528; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_530 = _instType_T_73 ? 5'h0 : _instType_T_529; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_531 = _instType_T_71 ? 5'h0 : _instType_T_530; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_532 = _instType_T_69 ? 5'h0 : _instType_T_531; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_533 = _instType_T_67 ? 5'h0 : _instType_T_532; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_534 = _instType_T_65 ? 5'h0 : _instType_T_533; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_535 = _instType_T_63 ? 5'h0 : _instType_T_534; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_536 = _instType_T_61 ? 5'h0 : _instType_T_535; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_537 = _instType_T_59 ? 5'h0 : _instType_T_536; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_538 = _instType_T_57 ? 5'h0 : _instType_T_537; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_539 = _instType_T_55 ? 5'h0 : _instType_T_538; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_540 = _instType_T_53 ? 5'h0 : _instType_T_539; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_541 = _instType_T_51 ? 5'h0 : _instType_T_540; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_542 = _instType_T_49 ? 5'h0 : _instType_T_541; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_543 = _instType_T_47 ? 5'h0 : _instType_T_542; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_544 = _instType_T_45 ? 5'h0 : _instType_T_543; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_545 = _instType_T_43 ? 5'h0 : _instType_T_544; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_546 = _instType_T_41 ? 5'hb : _instType_T_545; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_547 = _instType_T_39 ? 5'ha : _instType_T_546; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_548 = _instType_T_37 ? 5'h9 : _instType_T_547; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_549 = _instType_T_35 ? 5'h8 : _instType_T_548; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_550 = _instType_T_33 ? 5'h16 : _instType_T_549; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_551 = _instType_T_31 ? 5'h15 : _instType_T_550; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_552 = _instType_T_29 ? 5'h14 : _instType_T_551; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_553 = _instType_T_27 ? 5'h7 : _instType_T_552; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_554 = _instType_T_25 ? 5'h6 : _instType_T_553; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_555 = _instType_T_23 ? 5'h5 : _instType_T_554; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_556 = _instType_T_21 ? 5'h4 : _instType_T_555; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_557 = _instType_T_19 ? 5'h0 : _instType_T_556; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_558 = _instType_T_17 ? 5'h0 : _instType_T_557; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_559 = _instType_T_15 ? 5'h0 : _instType_T_558; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_560 = _instType_T_13 ? 5'h0 : _instType_T_559; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_561 = _instType_T_11 ? 5'h0 : _instType_T_560; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_562 = _instType_T_9 ? 5'h0 : _instType_T_561; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_563 = _instType_T_7 ? 5'h0 : _instType_T_562; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_564 = _instType_T_5 ? 5'h0 : _instType_T_563; // @[Lookup.scala 33:37]
  wire [4:0] _instType_T_565 = _instType_T_3 ? 5'h0 : _instType_T_564; // @[Lookup.scala 33:37]
  wire [4:0] instType_3 = _instType_T_1 ? 5'h0 : _instType_T_565; // @[Lookup.scala 33:37]
  wire  _instType_T_601 = _instType_T_119 | (_instType_T_121 | (_instType_T_123 | (_instType_T_125 | (_instType_T_127 |
    (_instType_T_129 | (_instType_T_131 | (_instType_T_133 | (_instType_T_135 | (_instType_T_137 | (_instType_T_139 | (
    _instType_T_141 | (_instType_T_143 | (_instType_T_145 | (_instType_T_147 | (_instType_T_149 | (_instType_T_151 | (
    _instType_T_153 | (_instType_T_155 | (_instType_T_157 | (_instType_T_159 | (_instType_T_161 | (_instType_T_163 | (
    _instType_T_165 | (_instType_T_167 | (_instType_T_169 | (_instType_T_171 | (_instType_T_173 | (_instType_T_175 | (
    _instType_T_177 | _instType_T_179))))))))))))))))))))))))))))); // @[Lookup.scala 33:37]
  wire  _instType_T_631 = _instType_T_59 | (_instType_T_61 | (_instType_T_63 | (_instType_T_65 | (_instType_T_67 | (
    _instType_T_69 | (_instType_T_71 | (_instType_T_73 | (_instType_T_75 | (_instType_T_77 | (_instType_T_79 | (
    _instType_T_81 | (_instType_T_83 | (_instType_T_85 | (_instType_T_87 | (_instType_T_89 | (_instType_T_91 | (
    _instType_T_93 | (_instType_T_95 | (_instType_T_97 | (_instType_T_99 | (_instType_T_101 | (_instType_T_103 | (
    _instType_T_105 | (_instType_T_107 | (_instType_T_109 | (_instType_T_111 | (_instType_T_113 | (_instType_T_115 | (
    _instType_T_117 | _instType_T_601))))))))))))))))))))))))))))); // @[Lookup.scala 33:37]
  wire  _instType_T_640 = _instType_T_41 ? 1'h0 : _instType_T_43 | (_instType_T_45 | (_instType_T_47 | (_instType_T_49
     | (_instType_T_51 | (_instType_T_53 | (_instType_T_55 | (_instType_T_57 | _instType_T_631))))))); // @[Lookup.scala 33:37]
  wire  _instType_T_641 = _instType_T_39 ? 1'h0 : _instType_T_640; // @[Lookup.scala 33:37]
  wire  _instType_T_642 = _instType_T_37 ? 1'h0 : _instType_T_641; // @[Lookup.scala 33:37]
  wire  _instType_T_643 = _instType_T_35 ? 1'h0 : _instType_T_642; // @[Lookup.scala 33:37]
  wire  _instType_T_651 = _instType_T_19 ? 1'h0 : _instType_T_21 | (_instType_T_23 | (_instType_T_25 | (_instType_T_27
     | (_instType_T_29 | (_instType_T_31 | (_instType_T_33 | _instType_T_643)))))); // @[Lookup.scala 33:37]
  wire  _instType_T_652 = _instType_T_17 ? 1'h0 : _instType_T_651; // @[Lookup.scala 33:37]
  wire  _instType_T_653 = _instType_T_15 ? 1'h0 : _instType_T_652; // @[Lookup.scala 33:37]
  wire  _instType_T_654 = _instType_T_13 ? 1'h0 : _instType_T_653; // @[Lookup.scala 33:37]
  wire  _instType_T_655 = _instType_T_11 ? 1'h0 : _instType_T_654; // @[Lookup.scala 33:37]
  wire  _instType_T_656 = _instType_T_9 ? 1'h0 : _instType_T_655; // @[Lookup.scala 33:37]
  wire  instType_4 = _instType_T_1 | (_instType_T_3 | (_instType_T_5 | (_instType_T_7 | _instType_T_656))); // @[Lookup.scala 33:37]
  wire  _instType_T_753 = _instType_T_3 ? 1'h0 : _instType_T_5 | (_instType_T_7 | (_instType_T_9 | (_instType_T_11 | (
    _instType_T_13 | (_instType_T_15 | (_instType_T_17 | _instType_T_19)))))); // @[Lookup.scala 33:37]
  wire  instType_5 = _instType_T_1 ? 1'h0 : _instType_T_753; // @[Lookup.scala 33:37]
  wire  _instType_T_787 = _instType_T_123 ? 1'h0 : _instType_T_125 | (_instType_T_127 | (_instType_T_129 | (
    _instType_T_131 | (_instType_T_133 | _instType_T_135)))); // @[Lookup.scala 33:37]
  wire  _instType_T_788 = _instType_T_121 ? 1'h0 : _instType_T_787; // @[Lookup.scala 33:37]
  wire  _instType_T_789 = _instType_T_119 ? 1'h0 : _instType_T_788; // @[Lookup.scala 33:37]
  wire  _instType_T_790 = _instType_T_117 ? 1'h0 : _instType_T_789; // @[Lookup.scala 33:37]
  wire  _instType_T_791 = _instType_T_115 ? 1'h0 : _instType_T_790; // @[Lookup.scala 33:37]
  wire  _instType_T_792 = _instType_T_113 ? 1'h0 : _instType_T_791; // @[Lookup.scala 33:37]
  wire  _instType_T_793 = _instType_T_111 ? 1'h0 : _instType_T_792; // @[Lookup.scala 33:37]
  wire  _instType_T_794 = _instType_T_109 ? 1'h0 : _instType_T_793; // @[Lookup.scala 33:37]
  wire  _instType_T_795 = _instType_T_107 ? 1'h0 : _instType_T_794; // @[Lookup.scala 33:37]
  wire  _instType_T_796 = _instType_T_105 ? 1'h0 : _instType_T_795; // @[Lookup.scala 33:37]
  wire  _instType_T_797 = _instType_T_103 ? 1'h0 : _instType_T_796; // @[Lookup.scala 33:37]
  wire  _instType_T_798 = _instType_T_101 ? 1'h0 : _instType_T_797; // @[Lookup.scala 33:37]
  wire  _instType_T_799 = _instType_T_99 ? 1'h0 : _instType_T_798; // @[Lookup.scala 33:37]
  wire  _instType_T_800 = _instType_T_97 ? 1'h0 : _instType_T_799; // @[Lookup.scala 33:37]
  wire  _instType_T_801 = _instType_T_95 ? 1'h0 : _instType_T_800; // @[Lookup.scala 33:37]
  wire  _instType_T_802 = _instType_T_93 ? 1'h0 : _instType_T_801; // @[Lookup.scala 33:37]
  wire  _instType_T_803 = _instType_T_91 ? 1'h0 : _instType_T_802; // @[Lookup.scala 33:37]
  wire  _instType_T_804 = _instType_T_89 ? 1'h0 : _instType_T_803; // @[Lookup.scala 33:37]
  wire  _instType_T_805 = _instType_T_87 ? 1'h0 : _instType_T_804; // @[Lookup.scala 33:37]
  wire  _instType_T_806 = _instType_T_85 ? 1'h0 : _instType_T_805; // @[Lookup.scala 33:37]
  wire  _instType_T_807 = _instType_T_83 ? 1'h0 : _instType_T_806; // @[Lookup.scala 33:37]
  wire  _instType_T_808 = _instType_T_81 ? 1'h0 : _instType_T_807; // @[Lookup.scala 33:37]
  wire  _instType_T_809 = _instType_T_79 ? 1'h0 : _instType_T_808; // @[Lookup.scala 33:37]
  wire  _instType_T_810 = _instType_T_77 ? 1'h0 : _instType_T_809; // @[Lookup.scala 33:37]
  wire  _instType_T_811 = _instType_T_75 ? 1'h0 : _instType_T_810; // @[Lookup.scala 33:37]
  wire  _instType_T_812 = _instType_T_73 ? 1'h0 : _instType_T_811; // @[Lookup.scala 33:37]
  wire  _instType_T_813 = _instType_T_71 ? 1'h0 : _instType_T_812; // @[Lookup.scala 33:37]
  wire  _instType_T_814 = _instType_T_69 ? 1'h0 : _instType_T_813; // @[Lookup.scala 33:37]
  wire  _instType_T_815 = _instType_T_67 ? 1'h0 : _instType_T_814; // @[Lookup.scala 33:37]
  wire  _instType_T_816 = _instType_T_65 ? 1'h0 : _instType_T_815; // @[Lookup.scala 33:37]
  wire  _instType_T_817 = _instType_T_63 ? 1'h0 : _instType_T_816; // @[Lookup.scala 33:37]
  wire  _instType_T_818 = _instType_T_61 ? 1'h0 : _instType_T_817; // @[Lookup.scala 33:37]
  wire  _instType_T_819 = _instType_T_59 ? 1'h0 : _instType_T_818; // @[Lookup.scala 33:37]
  wire  _instType_T_820 = _instType_T_57 ? 1'h0 : _instType_T_819; // @[Lookup.scala 33:37]
  wire  _instType_T_821 = _instType_T_55 ? 1'h0 : _instType_T_820; // @[Lookup.scala 33:37]
  wire  _instType_T_822 = _instType_T_53 ? 1'h0 : _instType_T_821; // @[Lookup.scala 33:37]
  wire  _instType_T_823 = _instType_T_51 ? 1'h0 : _instType_T_822; // @[Lookup.scala 33:37]
  wire  _instType_T_824 = _instType_T_49 ? 1'h0 : _instType_T_823; // @[Lookup.scala 33:37]
  wire  _instType_T_825 = _instType_T_47 ? 1'h0 : _instType_T_824; // @[Lookup.scala 33:37]
  wire  _instType_T_826 = _instType_T_45 ? 1'h0 : _instType_T_825; // @[Lookup.scala 33:37]
  wire  _instType_T_827 = _instType_T_43 ? 1'h0 : _instType_T_826; // @[Lookup.scala 33:37]
  wire  _instType_T_828 = _instType_T_41 ? 1'h0 : _instType_T_827; // @[Lookup.scala 33:37]
  wire  _instType_T_829 = _instType_T_39 ? 1'h0 : _instType_T_828; // @[Lookup.scala 33:37]
  wire  _instType_T_830 = _instType_T_37 ? 1'h0 : _instType_T_829; // @[Lookup.scala 33:37]
  wire  _instType_T_831 = _instType_T_35 ? 1'h0 : _instType_T_830; // @[Lookup.scala 33:37]
  wire  _instType_T_832 = _instType_T_33 ? 1'h0 : _instType_T_831; // @[Lookup.scala 33:37]
  wire  _instType_T_833 = _instType_T_31 ? 1'h0 : _instType_T_832; // @[Lookup.scala 33:37]
  wire  _instType_T_834 = _instType_T_29 ? 1'h0 : _instType_T_833; // @[Lookup.scala 33:37]
  wire  _instType_T_835 = _instType_T_27 ? 1'h0 : _instType_T_834; // @[Lookup.scala 33:37]
  wire  _instType_T_836 = _instType_T_25 ? 1'h0 : _instType_T_835; // @[Lookup.scala 33:37]
  wire  _instType_T_837 = _instType_T_23 ? 1'h0 : _instType_T_836; // @[Lookup.scala 33:37]
  wire  _instType_T_838 = _instType_T_21 ? 1'h0 : _instType_T_837; // @[Lookup.scala 33:37]
  wire  _instType_T_839 = _instType_T_19 ? 1'h0 : _instType_T_838; // @[Lookup.scala 33:37]
  wire  _instType_T_840 = _instType_T_17 ? 1'h0 : _instType_T_839; // @[Lookup.scala 33:37]
  wire  _instType_T_841 = _instType_T_15 ? 1'h0 : _instType_T_840; // @[Lookup.scala 33:37]
  wire  _instType_T_842 = _instType_T_13 ? 1'h0 : _instType_T_841; // @[Lookup.scala 33:37]
  wire  _instType_T_843 = _instType_T_11 ? 1'h0 : _instType_T_842; // @[Lookup.scala 33:37]
  wire  _instType_T_844 = _instType_T_9 ? 1'h0 : _instType_T_843; // @[Lookup.scala 33:37]
  wire  _instType_T_845 = _instType_T_7 ? 1'h0 : _instType_T_844; // @[Lookup.scala 33:37]
  wire  _instType_T_846 = _instType_T_5 ? 1'h0 : _instType_T_845; // @[Lookup.scala 33:37]
  wire  _instType_T_847 = _instType_T_3 ? 1'h0 : _instType_T_846; // @[Lookup.scala 33:37]
  wire  instType_6 = _instType_T_1 ? 1'h0 : _instType_T_847; // @[Lookup.scala 33:37]
  wire  _instType_T_972 = _instType_T_129 ? 1'h0 : _instType_T_131 | (_instType_T_133 | _instType_T_135); // @[Lookup.scala 33:37]
  wire  _instType_T_973 = _instType_T_127 ? 1'h0 : _instType_T_972; // @[Lookup.scala 33:37]
  wire  _instType_T_974 = _instType_T_125 ? 1'h0 : _instType_T_973; // @[Lookup.scala 33:37]
  wire  _instType_T_975 = _instType_T_123 ? 1'h0 : _instType_T_974; // @[Lookup.scala 33:37]
  wire  _instType_T_976 = _instType_T_121 ? 1'h0 : _instType_T_975; // @[Lookup.scala 33:37]
  wire  _instType_T_977 = _instType_T_119 ? 1'h0 : _instType_T_976; // @[Lookup.scala 33:37]
  wire  _instType_T_978 = _instType_T_117 ? 1'h0 : _instType_T_977; // @[Lookup.scala 33:37]
  wire  _instType_T_979 = _instType_T_115 ? 1'h0 : _instType_T_978; // @[Lookup.scala 33:37]
  wire  _instType_T_980 = _instType_T_113 ? 1'h0 : _instType_T_979; // @[Lookup.scala 33:37]
  wire  _instType_T_981 = _instType_T_111 ? 1'h0 : _instType_T_980; // @[Lookup.scala 33:37]
  wire  _instType_T_982 = _instType_T_109 ? 1'h0 : _instType_T_981; // @[Lookup.scala 33:37]
  wire  _instType_T_983 = _instType_T_107 ? 1'h0 : _instType_T_982; // @[Lookup.scala 33:37]
  wire  _instType_T_984 = _instType_T_105 ? 1'h0 : _instType_T_983; // @[Lookup.scala 33:37]
  wire  _instType_T_985 = _instType_T_103 ? 1'h0 : _instType_T_984; // @[Lookup.scala 33:37]
  wire  _instType_T_986 = _instType_T_101 ? 1'h0 : _instType_T_985; // @[Lookup.scala 33:37]
  wire  _instType_T_987 = _instType_T_99 ? 1'h0 : _instType_T_986; // @[Lookup.scala 33:37]
  wire  _instType_T_988 = _instType_T_97 ? 1'h0 : _instType_T_987; // @[Lookup.scala 33:37]
  wire  _instType_T_989 = _instType_T_95 ? 1'h0 : _instType_T_988; // @[Lookup.scala 33:37]
  wire  _instType_T_990 = _instType_T_93 ? 1'h0 : _instType_T_989; // @[Lookup.scala 33:37]
  wire  _instType_T_991 = _instType_T_91 ? 1'h0 : _instType_T_990; // @[Lookup.scala 33:37]
  wire  _instType_T_992 = _instType_T_89 ? 1'h0 : _instType_T_991; // @[Lookup.scala 33:37]
  wire  _instType_T_993 = _instType_T_87 ? 1'h0 : _instType_T_992; // @[Lookup.scala 33:37]
  wire  _instType_T_994 = _instType_T_85 ? 1'h0 : _instType_T_993; // @[Lookup.scala 33:37]
  wire  _instType_T_995 = _instType_T_83 ? 1'h0 : _instType_T_994; // @[Lookup.scala 33:37]
  wire  _instType_T_996 = _instType_T_81 ? 1'h0 : _instType_T_995; // @[Lookup.scala 33:37]
  wire  _instType_T_997 = _instType_T_79 ? 1'h0 : _instType_T_996; // @[Lookup.scala 33:37]
  wire  _instType_T_998 = _instType_T_77 ? 1'h0 : _instType_T_997; // @[Lookup.scala 33:37]
  wire  _instType_T_999 = _instType_T_75 ? 1'h0 : _instType_T_998; // @[Lookup.scala 33:37]
  wire  _instType_T_1000 = _instType_T_73 ? 1'h0 : _instType_T_999; // @[Lookup.scala 33:37]
  wire  _instType_T_1001 = _instType_T_71 ? 1'h0 : _instType_T_1000; // @[Lookup.scala 33:37]
  wire  _instType_T_1002 = _instType_T_69 ? 1'h0 : _instType_T_1001; // @[Lookup.scala 33:37]
  wire  _instType_T_1003 = _instType_T_67 ? 1'h0 : _instType_T_1002; // @[Lookup.scala 33:37]
  wire  _instType_T_1004 = _instType_T_65 ? 1'h0 : _instType_T_1003; // @[Lookup.scala 33:37]
  wire  _instType_T_1005 = _instType_T_63 ? 1'h0 : _instType_T_1004; // @[Lookup.scala 33:37]
  wire  _instType_T_1006 = _instType_T_61 ? 1'h0 : _instType_T_1005; // @[Lookup.scala 33:37]
  wire  _instType_T_1007 = _instType_T_59 ? 1'h0 : _instType_T_1006; // @[Lookup.scala 33:37]
  wire  _instType_T_1008 = _instType_T_57 ? 1'h0 : _instType_T_1007; // @[Lookup.scala 33:37]
  wire  _instType_T_1009 = _instType_T_55 ? 1'h0 : _instType_T_1008; // @[Lookup.scala 33:37]
  wire  _instType_T_1010 = _instType_T_53 ? 1'h0 : _instType_T_1009; // @[Lookup.scala 33:37]
  wire  _instType_T_1011 = _instType_T_51 ? 1'h0 : _instType_T_1010; // @[Lookup.scala 33:37]
  wire  _instType_T_1012 = _instType_T_49 ? 1'h0 : _instType_T_1011; // @[Lookup.scala 33:37]
  wire  _instType_T_1013 = _instType_T_47 ? 1'h0 : _instType_T_1012; // @[Lookup.scala 33:37]
  wire  _instType_T_1014 = _instType_T_45 ? 1'h0 : _instType_T_1013; // @[Lookup.scala 33:37]
  wire  _instType_T_1015 = _instType_T_43 ? 1'h0 : _instType_T_1014; // @[Lookup.scala 33:37]
  wire  _instType_T_1016 = _instType_T_41 ? 1'h0 : _instType_T_1015; // @[Lookup.scala 33:37]
  wire  _instType_T_1017 = _instType_T_39 ? 1'h0 : _instType_T_1016; // @[Lookup.scala 33:37]
  wire  _instType_T_1018 = _instType_T_37 ? 1'h0 : _instType_T_1017; // @[Lookup.scala 33:37]
  wire  _instType_T_1019 = _instType_T_35 ? 1'h0 : _instType_T_1018; // @[Lookup.scala 33:37]
  wire  _instType_T_1020 = _instType_T_33 ? 1'h0 : _instType_T_1019; // @[Lookup.scala 33:37]
  wire  _instType_T_1021 = _instType_T_31 ? 1'h0 : _instType_T_1020; // @[Lookup.scala 33:37]
  wire  _instType_T_1022 = _instType_T_29 ? 1'h0 : _instType_T_1021; // @[Lookup.scala 33:37]
  wire  _instType_T_1023 = _instType_T_27 ? 1'h0 : _instType_T_1022; // @[Lookup.scala 33:37]
  wire  _instType_T_1024 = _instType_T_25 ? 1'h0 : _instType_T_1023; // @[Lookup.scala 33:37]
  wire  _instType_T_1025 = _instType_T_23 ? 1'h0 : _instType_T_1024; // @[Lookup.scala 33:37]
  wire  _instType_T_1026 = _instType_T_21 ? 1'h0 : _instType_T_1025; // @[Lookup.scala 33:37]
  wire  _instType_T_1027 = _instType_T_19 ? 1'h0 : _instType_T_1026; // @[Lookup.scala 33:37]
  wire  _instType_T_1028 = _instType_T_17 ? 1'h0 : _instType_T_1027; // @[Lookup.scala 33:37]
  wire  _instType_T_1029 = _instType_T_15 ? 1'h0 : _instType_T_1028; // @[Lookup.scala 33:37]
  wire  _instType_T_1030 = _instType_T_13 ? 1'h0 : _instType_T_1029; // @[Lookup.scala 33:37]
  wire  _instType_T_1031 = _instType_T_11 ? 1'h0 : _instType_T_1030; // @[Lookup.scala 33:37]
  wire  _instType_T_1032 = _instType_T_9 ? 1'h0 : _instType_T_1031; // @[Lookup.scala 33:37]
  wire  _instType_T_1033 = _instType_T_7 ? 1'h0 : _instType_T_1032; // @[Lookup.scala 33:37]
  wire  _instType_T_1034 = _instType_T_5 ? 1'h0 : _instType_T_1033; // @[Lookup.scala 33:37]
  wire  _instType_T_1035 = _instType_T_3 ? 1'h0 : _instType_T_1034; // @[Lookup.scala 33:37]
  wire  instType_8 = _instType_T_1 ? 1'h0 : _instType_T_1035; // @[Lookup.scala 33:37]
  wire [15:0] _instType_c_T_1 = io_if2id_inst[15:0] & 16'he003; // @[Lookup.scala 31:38]
  wire  _instType_c_T_2 = 16'h0 == _instType_c_T_1; // @[Lookup.scala 31:38]
  wire  _instType_c_T_4 = 16'h4000 == _instType_c_T_1; // @[Lookup.scala 31:38]
  wire  _instType_c_T_6 = 16'h6000 == _instType_c_T_1; // @[Lookup.scala 31:38]
  wire  _instType_c_T_8 = 16'hc000 == _instType_c_T_1; // @[Lookup.scala 31:38]
  wire  _instType_c_T_10 = 16'he000 == _instType_c_T_1; // @[Lookup.scala 31:38]
  wire  _instType_c_T_12 = 16'h1 == _instType_c_T_1; // @[Lookup.scala 31:38]
  wire  _instType_c_T_14 = 16'h2001 == _instType_c_T_1; // @[Lookup.scala 31:38]
  wire  _instType_c_T_16 = 16'h4001 == _instType_c_T_1; // @[Lookup.scala 31:38]
  wire [15:0] _instType_c_T_17 = io_if2id_inst[15:0] & 16'hef83; // @[Lookup.scala 31:38]
  wire  _instType_c_T_18 = 16'h6101 == _instType_c_T_17; // @[Lookup.scala 31:38]
  wire  _instType_c_T_20 = 16'h6001 == _instType_c_T_1; // @[Lookup.scala 31:38]
  wire [15:0] _instType_c_T_21 = io_if2id_inst[15:0] & 16'hec03; // @[Lookup.scala 31:38]
  wire  _instType_c_T_22 = 16'h8001 == _instType_c_T_21; // @[Lookup.scala 31:38]
  wire  _instType_c_T_24 = 16'h8401 == _instType_c_T_21; // @[Lookup.scala 31:38]
  wire  _instType_c_T_26 = 16'h8801 == _instType_c_T_21; // @[Lookup.scala 31:38]
  wire [15:0] _instType_c_T_27 = io_if2id_inst[15:0] & 16'hfc63; // @[Lookup.scala 31:38]
  wire  _instType_c_T_28 = 16'h8c01 == _instType_c_T_27; // @[Lookup.scala 31:38]
  wire  _instType_c_T_30 = 16'h8c21 == _instType_c_T_27; // @[Lookup.scala 31:38]
  wire  _instType_c_T_32 = 16'h8c41 == _instType_c_T_27; // @[Lookup.scala 31:38]
  wire  _instType_c_T_34 = 16'h8c61 == _instType_c_T_27; // @[Lookup.scala 31:38]
  wire  _instType_c_T_36 = 16'h9c01 == _instType_c_T_27; // @[Lookup.scala 31:38]
  wire  _instType_c_T_38 = 16'h9c21 == _instType_c_T_27; // @[Lookup.scala 31:38]
  wire  _instType_c_T_40 = 16'ha001 == _instType_c_T_1; // @[Lookup.scala 31:38]
  wire  _instType_c_T_42 = 16'hc001 == _instType_c_T_1; // @[Lookup.scala 31:38]
  wire  _instType_c_T_44 = 16'he001 == _instType_c_T_1; // @[Lookup.scala 31:38]
  wire  _instType_c_T_46 = 16'h2 == _instType_c_T_1; // @[Lookup.scala 31:38]
  wire  _instType_c_T_48 = 16'h4002 == _instType_c_T_1; // @[Lookup.scala 31:38]
  wire  _instType_c_T_50 = 16'h6002 == _instType_c_T_1; // @[Lookup.scala 31:38]
  wire [15:0] _instType_c_T_51 = io_if2id_inst[15:0] & 16'hf07f; // @[Lookup.scala 31:38]
  wire  _instType_c_T_52 = 16'h8002 == _instType_c_T_51; // @[Lookup.scala 31:38]
  wire [15:0] _instType_c_T_53 = io_if2id_inst[15:0] & 16'hf003; // @[Lookup.scala 31:38]
  wire  _instType_c_T_54 = 16'h8002 == _instType_c_T_53; // @[Lookup.scala 31:38]
  wire  _instType_c_T_56 = 16'h9002 == _instType_c_T_51; // @[Lookup.scala 31:38]
  wire  _instType_c_T_58 = 16'h9002 == _instType_c_T_53; // @[Lookup.scala 31:38]
  wire  _instType_c_T_60 = 16'hc002 == _instType_c_T_1; // @[Lookup.scala 31:38]
  wire  _instType_c_T_62 = 16'he002 == _instType_c_T_1; // @[Lookup.scala 31:38]
  wire [3:0] _instType_c_T_63 = _instType_c_T_62 ? 4'h3 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_64 = _instType_c_T_60 ? 4'h3 : _instType_c_T_63; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_65 = _instType_c_T_58 ? 4'h1 : _instType_c_T_64; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_66 = _instType_c_T_56 ? 4'h1 : _instType_c_T_65; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_67 = _instType_c_T_54 ? 4'h1 : _instType_c_T_66; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_68 = _instType_c_T_52 ? 4'h1 : _instType_c_T_67; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_69 = _instType_c_T_50 ? 4'h2 : _instType_c_T_68; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_70 = _instType_c_T_48 ? 4'h2 : _instType_c_T_69; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_71 = _instType_c_T_46 ? 4'h2 : _instType_c_T_70; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_72 = _instType_c_T_44 ? 4'h7 : _instType_c_T_71; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_73 = _instType_c_T_42 ? 4'h7 : _instType_c_T_72; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_74 = _instType_c_T_40 ? 4'h8 : _instType_c_T_73; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_75 = _instType_c_T_38 ? 4'h6 : _instType_c_T_74; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_76 = _instType_c_T_36 ? 4'h6 : _instType_c_T_75; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_77 = _instType_c_T_34 ? 4'h6 : _instType_c_T_76; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_78 = _instType_c_T_32 ? 4'h6 : _instType_c_T_77; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_79 = _instType_c_T_30 ? 4'h6 : _instType_c_T_78; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_80 = _instType_c_T_28 ? 4'h6 : _instType_c_T_79; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_81 = _instType_c_T_26 ? 4'h7 : _instType_c_T_80; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_82 = _instType_c_T_24 ? 4'h7 : _instType_c_T_81; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_83 = _instType_c_T_22 ? 4'h7 : _instType_c_T_82; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_84 = _instType_c_T_20 ? 4'h2 : _instType_c_T_83; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_85 = _instType_c_T_18 ? 4'h2 : _instType_c_T_84; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_86 = _instType_c_T_16 ? 4'h2 : _instType_c_T_85; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_87 = _instType_c_T_14 ? 4'h2 : _instType_c_T_86; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_88 = _instType_c_T_12 ? 4'h2 : _instType_c_T_87; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_89 = _instType_c_T_10 ? 4'h6 : _instType_c_T_88; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_90 = _instType_c_T_8 ? 4'h6 : _instType_c_T_89; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_91 = _instType_c_T_6 ? 4'h5 : _instType_c_T_90; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_92 = _instType_c_T_4 ? 4'h5 : _instType_c_T_91; // @[Lookup.scala 33:37]
  wire [3:0] instType_c_0 = _instType_c_T_2 ? 4'h4 : _instType_c_T_92; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_93 = _instType_c_T_62 ? 4'hd : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_94 = _instType_c_T_60 ? 4'hc : _instType_c_T_93; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_95 = _instType_c_T_58 ? 4'h0 : _instType_c_T_94; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_96 = _instType_c_T_56 ? 4'h0 : _instType_c_T_95; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_97 = _instType_c_T_54 ? 4'h0 : _instType_c_T_96; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_98 = _instType_c_T_52 ? 4'h0 : _instType_c_T_97; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_99 = _instType_c_T_50 ? 4'h7 : _instType_c_T_98; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_100 = _instType_c_T_48 ? 4'h6 : _instType_c_T_99; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_101 = _instType_c_T_46 ? 4'h4 : _instType_c_T_100; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_102 = _instType_c_T_44 ? 4'hb : _instType_c_T_101; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_103 = _instType_c_T_42 ? 4'hb : _instType_c_T_102; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_104 = _instType_c_T_40 ? 4'ha : _instType_c_T_103; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_105 = _instType_c_T_38 ? 4'h0 : _instType_c_T_104; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_106 = _instType_c_T_36 ? 4'h0 : _instType_c_T_105; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_107 = _instType_c_T_34 ? 4'h0 : _instType_c_T_106; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_108 = _instType_c_T_32 ? 4'h0 : _instType_c_T_107; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_109 = _instType_c_T_30 ? 4'h0 : _instType_c_T_108; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_110 = _instType_c_T_28 ? 4'h0 : _instType_c_T_109; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_111 = _instType_c_T_26 ? 4'h5 : _instType_c_T_110; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_112 = _instType_c_T_24 ? 4'h4 : _instType_c_T_111; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_113 = _instType_c_T_22 ? 4'h4 : _instType_c_T_112; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_114 = _instType_c_T_20 ? 4'h9 : _instType_c_T_113; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_115 = _instType_c_T_18 ? 4'h8 : _instType_c_T_114; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_116 = _instType_c_T_16 ? 4'h5 : _instType_c_T_115; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_117 = _instType_c_T_14 ? 4'h5 : _instType_c_T_116; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_118 = _instType_c_T_12 ? 4'h5 : _instType_c_T_117; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_119 = _instType_c_T_10 ? 4'h3 : _instType_c_T_118; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_120 = _instType_c_T_8 ? 4'h2 : _instType_c_T_119; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_121 = _instType_c_T_6 ? 4'h3 : _instType_c_T_120; // @[Lookup.scala 33:37]
  wire [3:0] _instType_c_T_122 = _instType_c_T_4 ? 4'h2 : _instType_c_T_121; // @[Lookup.scala 33:37]
  wire [3:0] instType_c_1 = _instType_c_T_2 ? 4'h1 : _instType_c_T_122; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_123 = _instType_c_T_62 ? 5'h3 : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_124 = _instType_c_T_60 ? 5'h3 : _instType_c_T_123; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_125 = _instType_c_T_58 ? 5'h3 : _instType_c_T_124; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_126 = _instType_c_T_56 ? 5'h2 : _instType_c_T_125; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_127 = _instType_c_T_54 ? 5'h2 : _instType_c_T_126; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_128 = _instType_c_T_52 ? 5'h1 : _instType_c_T_127; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_129 = _instType_c_T_50 ? 5'h3 : _instType_c_T_128; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_130 = _instType_c_T_48 ? 5'h3 : _instType_c_T_129; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_131 = _instType_c_T_46 ? 5'h7 : _instType_c_T_130; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_132 = _instType_c_T_44 ? 5'h0 : _instType_c_T_131; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_133 = _instType_c_T_42 ? 5'h0 : _instType_c_T_132; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_134 = _instType_c_T_40 ? 5'h2 : _instType_c_T_133; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_135 = _instType_c_T_38 ? 5'h3 : _instType_c_T_134; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_136 = _instType_c_T_36 ? 5'ha : _instType_c_T_135; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_137 = _instType_c_T_34 ? 5'h6 : _instType_c_T_136; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_138 = _instType_c_T_32 ? 5'h5 : _instType_c_T_137; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_139 = _instType_c_T_30 ? 5'h4 : _instType_c_T_138; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_140 = _instType_c_T_28 ? 5'ha : _instType_c_T_139; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_141 = _instType_c_T_26 ? 5'h6 : _instType_c_T_140; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_142 = _instType_c_T_24 ? 5'h9 : _instType_c_T_141; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_143 = _instType_c_T_22 ? 5'h8 : _instType_c_T_142; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_144 = _instType_c_T_20 ? 5'h2 : _instType_c_T_143; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_145 = _instType_c_T_18 ? 5'h3 : _instType_c_T_144; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_146 = _instType_c_T_16 ? 5'h2 : _instType_c_T_145; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_147 = _instType_c_T_14 ? 5'h3 : _instType_c_T_146; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_148 = _instType_c_T_12 ? 5'h3 : _instType_c_T_147; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_149 = _instType_c_T_10 ? 5'h3 : _instType_c_T_148; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_150 = _instType_c_T_8 ? 5'h3 : _instType_c_T_149; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_151 = _instType_c_T_6 ? 5'h3 : _instType_c_T_150; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_152 = _instType_c_T_4 ? 5'h3 : _instType_c_T_151; // @[Lookup.scala 33:37]
  wire  _instType_c_T_167 = _instType_c_T_34 ? 1'h0 : _instType_c_T_36 | _instType_c_T_38; // @[Lookup.scala 33:37]
  wire  _instType_c_T_168 = _instType_c_T_32 ? 1'h0 : _instType_c_T_167; // @[Lookup.scala 33:37]
  wire  _instType_c_T_169 = _instType_c_T_30 ? 1'h0 : _instType_c_T_168; // @[Lookup.scala 33:37]
  wire  _instType_c_T_170 = _instType_c_T_28 ? 1'h0 : _instType_c_T_169; // @[Lookup.scala 33:37]
  wire  _instType_c_T_171 = _instType_c_T_26 ? 1'h0 : _instType_c_T_170; // @[Lookup.scala 33:37]
  wire  _instType_c_T_172 = _instType_c_T_24 ? 1'h0 : _instType_c_T_171; // @[Lookup.scala 33:37]
  wire  _instType_c_T_173 = _instType_c_T_22 ? 1'h0 : _instType_c_T_172; // @[Lookup.scala 33:37]
  wire  _instType_c_T_174 = _instType_c_T_20 ? 1'h0 : _instType_c_T_173; // @[Lookup.scala 33:37]
  wire  _instType_c_T_175 = _instType_c_T_18 ? 1'h0 : _instType_c_T_174; // @[Lookup.scala 33:37]
  wire  _instType_c_T_176 = _instType_c_T_16 ? 1'h0 : _instType_c_T_175; // @[Lookup.scala 33:37]
  wire  _instType_c_T_178 = _instType_c_T_12 ? 1'h0 : _instType_c_T_14 | _instType_c_T_176; // @[Lookup.scala 33:37]
  wire  _instType_c_T_179 = _instType_c_T_10 ? 1'h0 : _instType_c_T_178; // @[Lookup.scala 33:37]
  wire  _instType_c_T_180 = _instType_c_T_8 ? 1'h0 : _instType_c_T_179; // @[Lookup.scala 33:37]
  wire  _instType_c_T_181 = _instType_c_T_6 ? 1'h0 : _instType_c_T_180; // @[Lookup.scala 33:37]
  wire  _instType_c_T_182 = _instType_c_T_4 ? 1'h0 : _instType_c_T_181; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_183 = _instType_c_T_62 ? 5'hb : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_184 = _instType_c_T_60 ? 5'ha : _instType_c_T_183; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_185 = _instType_c_T_58 ? 5'h0 : _instType_c_T_184; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_186 = _instType_c_T_56 ? 5'h0 : _instType_c_T_185; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_187 = _instType_c_T_54 ? 5'h0 : _instType_c_T_186; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_188 = _instType_c_T_52 ? 5'h0 : _instType_c_T_187; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_189 = _instType_c_T_50 ? 5'h7 : _instType_c_T_188; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_190 = _instType_c_T_48 ? 5'h6 : _instType_c_T_189; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_191 = _instType_c_T_46 ? 5'h0 : _instType_c_T_190; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_192 = _instType_c_T_44 ? 5'h0 : _instType_c_T_191; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_193 = _instType_c_T_42 ? 5'h0 : _instType_c_T_192; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_194 = _instType_c_T_40 ? 5'h0 : _instType_c_T_193; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_195 = _instType_c_T_38 ? 5'h0 : _instType_c_T_194; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_196 = _instType_c_T_36 ? 5'h0 : _instType_c_T_195; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_197 = _instType_c_T_34 ? 5'h0 : _instType_c_T_196; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_198 = _instType_c_T_32 ? 5'h0 : _instType_c_T_197; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_199 = _instType_c_T_30 ? 5'h0 : _instType_c_T_198; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_200 = _instType_c_T_28 ? 5'h0 : _instType_c_T_199; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_201 = _instType_c_T_26 ? 5'h0 : _instType_c_T_200; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_202 = _instType_c_T_24 ? 5'h0 : _instType_c_T_201; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_203 = _instType_c_T_22 ? 5'h0 : _instType_c_T_202; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_204 = _instType_c_T_20 ? 5'h0 : _instType_c_T_203; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_205 = _instType_c_T_18 ? 5'h0 : _instType_c_T_204; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_206 = _instType_c_T_16 ? 5'h0 : _instType_c_T_205; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_207 = _instType_c_T_14 ? 5'h0 : _instType_c_T_206; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_208 = _instType_c_T_12 ? 5'h0 : _instType_c_T_207; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_209 = _instType_c_T_10 ? 5'hb : _instType_c_T_208; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_210 = _instType_c_T_8 ? 5'ha : _instType_c_T_209; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_211 = _instType_c_T_6 ? 5'h7 : _instType_c_T_210; // @[Lookup.scala 33:37]
  wire [4:0] _instType_c_T_212 = _instType_c_T_4 ? 5'h6 : _instType_c_T_211; // @[Lookup.scala 33:37]
  wire  _instType_c_T_218 = _instType_c_T_52 ? 1'h0 : _instType_c_T_54 | (_instType_c_T_56 | _instType_c_T_58); // @[Lookup.scala 33:37]
  wire  _instType_c_T_222 = _instType_c_T_44 ? 1'h0 : _instType_c_T_46 | (_instType_c_T_48 | (_instType_c_T_50 |
    _instType_c_T_218)); // @[Lookup.scala 33:37]
  wire  _instType_c_T_223 = _instType_c_T_42 ? 1'h0 : _instType_c_T_222; // @[Lookup.scala 33:37]
  wire  _instType_c_T_224 = _instType_c_T_40 ? 1'h0 : _instType_c_T_223; // @[Lookup.scala 33:37]
  wire  _instType_c_T_239 = _instType_c_T_10 ? 1'h0 : _instType_c_T_12 | (_instType_c_T_14 | (_instType_c_T_16 | (
    _instType_c_T_18 | (_instType_c_T_20 | (_instType_c_T_22 | (_instType_c_T_24 | (_instType_c_T_26 | (_instType_c_T_28
     | (_instType_c_T_30 | (_instType_c_T_32 | (_instType_c_T_34 | (_instType_c_T_36 | (_instType_c_T_38 |
    _instType_c_T_224))))))))))))); // @[Lookup.scala 33:37]
  wire  _instType_c_T_240 = _instType_c_T_8 ? 1'h0 : _instType_c_T_239; // @[Lookup.scala 33:37]
  wire  instType_c_5 = _instType_c_T_2 | (_instType_c_T_4 | (_instType_c_T_6 | _instType_c_T_240)); // @[Lookup.scala 33:37]
  wire  is_compress = io_if2id_inst[1:0] != 2'h3; // @[decode.scala 56:36]
  wire  _T = 3'h2 == dType; // @[Conditional.scala 37:30]
  wire [11:0] _imm_T_1 = io_if2id_inst[31:20]; // @[decode.scala 59:42]
  wire  _T_1 = 3'h3 == dType; // @[Conditional.scala 37:30]
  wire [6:0] imm_hi = io_if2id_inst[31:25]; // @[decode.scala 60:38]
  wire [4:0] imm_lo = io_if2id_inst[11:7]; // @[decode.scala 60:55]
  wire [11:0] _imm_T_3 = {imm_hi,imm_lo}; // @[decode.scala 60:64]
  wire  _T_2 = 3'h4 == dType; // @[Conditional.scala 37:30]
  wire  imm_hi_hi_hi = io_if2id_inst[31]; // @[decode.scala 61:38]
  wire  imm_hi_hi_lo = io_if2id_inst[7]; // @[decode.scala 61:51]
  wire [5:0] imm_hi_lo = io_if2id_inst[30:25]; // @[decode.scala 61:63]
  wire [3:0] imm_lo_hi = io_if2id_inst[11:8]; // @[decode.scala 61:80]
  wire [12:0] _imm_T_5 = {imm_hi_hi_hi,imm_hi_hi_lo,imm_hi_lo,imm_lo_hi,1'h0}; // @[decode.scala 61:99]
  wire  _T_3 = 3'h5 == dType; // @[Conditional.scala 37:30]
  wire [19:0] imm_hi_2 = io_if2id_inst[31:12]; // @[decode.scala 62:38]
  wire [31:0] _imm_T_7 = {imm_hi_2,12'h0}; // @[decode.scala 62:59]
  wire  _T_4 = 3'h6 == dType; // @[Conditional.scala 37:30]
  wire [7:0] imm_hi_hi_lo_1 = io_if2id_inst[19:12]; // @[decode.scala 63:51]
  wire  imm_hi_lo_1 = io_if2id_inst[20]; // @[decode.scala 63:68]
  wire [9:0] imm_lo_hi_1 = io_if2id_inst[30:21]; // @[decode.scala 63:81]
  wire [20:0] _imm_T_9 = {imm_hi_hi_hi,imm_hi_hi_lo_1,imm_hi_lo_1,imm_lo_hi_1,1'h0}; // @[decode.scala 63:101]
  wire [20:0] _GEN_0 = _T_4 ? $signed(_imm_T_9) : $signed(21'sh0); // @[Conditional.scala 39:67 decode.scala 63:24 decode.scala 57:9]
  wire [31:0] _GEN_1 = _T_3 ? $signed(_imm_T_7) : $signed({{11{_GEN_0[20]}},_GEN_0}); // @[Conditional.scala 39:67 decode.scala 62:24]
  wire [31:0] _GEN_2 = _T_2 ? $signed({{19{_imm_T_5[12]}},_imm_T_5}) : $signed(_GEN_1); // @[Conditional.scala 39:67 decode.scala 61:24]
  wire [31:0] _GEN_3 = _T_1 ? $signed({{20{_imm_T_3[11]}},_imm_T_3}) : $signed(_GEN_2); // @[Conditional.scala 39:67 decode.scala 60:24]
  wire [31:0] _GEN_4 = _T ? $signed({{20{_imm_T_1[11]}},_imm_T_1}) : $signed(_GEN_3); // @[Conditional.scala 40:58 decode.scala 59:24]
  wire  _T_7 = ~io_if2id_excep_en; // @[decode.scala 65:35]
  wire [11:0] _rs2_r_T_2 = instType_6 ? io_if2id_inst[31:20] : {{7'd0}, io_if2id_inst[24:20]}; // @[decode.scala 76:31]
  wire  indi_r_hi = _instType_T_139 | _instType_T_161; // @[decode.scala 81:55]
  wire  indi_r_lo = _instType_T_137 | _instType_T_159; // @[decode.scala 82:56]
  wire [1:0] _indi_r_T_8 = {indi_r_hi,indi_r_lo}; // @[Cat.scala 30:58]
  wire  _T_11 = dType == 3'h7 & _T_7; // @[decode.scala 85:32]
  wire  _GEN_5 = dType == 3'h7 & _T_7 | io_if2id_excep_en; // @[decode.scala 85:54 decode.scala 86:29 decode.scala 68:25]
  wire [63:0] _GEN_6 = dType == 3'h7 & _T_7 ? 64'h2 : io_if2id_excep_cause; // @[decode.scala 85:54 decode.scala 87:29 decode.scala 68:25]
  wire [63:0] _GEN_7 = dType == 3'h7 & _T_7 ? {{32'd0}, io_if2id_inst} : io_if2id_excep_tval; // @[decode.scala 85:54 decode.scala 88:29 decode.scala 68:25]
  wire [63:0] _GEN_8 = dType == 3'h7 & _T_7 ? io_if2id_pc : io_if2id_excep_pc; // @[decode.scala 85:54 decode.scala 89:29 decode.scala 68:25]
  wire  _GEN_11 = dType == 3'h7 & _T_7 | io_if2id_recov; // @[decode.scala 85:54 decode.scala 43:57 decode.scala 84:25]
  wire  _T_12 = dType == 3'h1; // @[decode.scala 93:20]
  wire [5:0] _GEN_13 = dType == 3'h1 ? 6'h1a : 6'h1b; // @[decode.scala 93:30 decode.scala 96:21 decode.scala 83:25]
  wire [63:0] _rs2_d_r_T_1 = io_if2id_pc + 64'h4; // @[decode.scala 102:44]
  wire [63:0] imm = {{32{_GEN_4[31]}},_GEN_4}; // @[decode.scala 55:19]
  wire [63:0] _dst_d_r_T = {{32{_GEN_4[31]}},_GEN_4}; // @[decode.scala 103:36]
  wire [63:0] _GEN_14 = instType_6 ? {{59'd0}, io_if2id_inst[19:15]} : rs1_d_r; // @[decode.scala 104:35 decode.scala 105:29 decode.scala 29:30]
  wire  _GEN_15 = instType_6 ? ~instType_8 : 1'h1; // @[decode.scala 104:35 decode.scala 106:29 decode.scala 110:29]
  wire  _GEN_16 = instType_6 | _T_12; // @[decode.scala 104:35 decode.scala 107:29]
  wire  _GEN_17 = instType_6 | _T_11; // @[decode.scala 104:35 decode.scala 43:17]
  wire  _GEN_18 = instType_6 | _GEN_11; // @[decode.scala 104:35 decode.scala 43:57]
  wire [63:0] _GEN_19 = instType_6 ? rs2_d_r : _dst_d_r_T; // @[decode.scala 104:35 decode.scala 32:30 decode.scala 111:29]
  wire [1:0] _GEN_20 = instType_5 ? 2'h1 : 2'h0; // @[decode.scala 99:27 decode.scala 100:29 decode.scala 79:25]
  wire  _GEN_21 = instType_5 | _GEN_15; // @[decode.scala 99:27 decode.scala 101:29]
  wire [63:0] _GEN_22 = instType_5 ? _rs2_d_r_T_1 : _GEN_19; // @[decode.scala 99:27 decode.scala 102:29]
  wire [63:0] _GEN_23 = instType_5 ? _dst_d_r_T : dst_d_r; // @[decode.scala 99:27 decode.scala 103:29 decode.scala 34:30]
  wire [63:0] _GEN_24 = instType_5 ? rs1_d_r : _GEN_14; // @[decode.scala 99:27 decode.scala 29:30]
  wire  _GEN_25 = instType_5 ? _T_12 : _GEN_16; // @[decode.scala 99:27]
  wire  _GEN_26 = instType_5 ? _T_11 : _GEN_17; // @[decode.scala 99:27]
  wire  _GEN_27 = instType_5 ? _GEN_11 : _GEN_18; // @[decode.scala 99:27]
  wire [1:0] _GEN_28 = dType == 3'h2 ? _GEN_20 : 2'h0; // @[decode.scala 98:30 decode.scala 79:25]
  wire  _GEN_29 = dType == 3'h2 ? _GEN_21 : _T_12; // @[decode.scala 98:30]
  wire [63:0] _GEN_30 = dType == 3'h2 ? _GEN_22 : rs2_d_r; // @[decode.scala 98:30 decode.scala 32:30]
  wire [63:0] _GEN_31 = dType == 3'h2 ? _GEN_23 : dst_d_r; // @[decode.scala 98:30 decode.scala 34:30]
  wire [63:0] _GEN_32 = dType == 3'h2 ? _GEN_24 : rs1_d_r; // @[decode.scala 98:30 decode.scala 29:30]
  wire  _GEN_33 = dType == 3'h2 ? _GEN_25 : _T_12; // @[decode.scala 98:30]
  wire  _GEN_34 = dType == 3'h2 ? _GEN_26 : _T_11; // @[decode.scala 98:30]
  wire  _GEN_35 = dType == 3'h2 ? _GEN_27 : _GEN_11; // @[decode.scala 98:30]
  wire  _GEN_36 = dType == 3'h3 | _GEN_29; // @[decode.scala 114:30 decode.scala 115:25]
  wire  _GEN_37 = dType == 3'h3 | _GEN_33; // @[decode.scala 114:30 decode.scala 116:25]
  wire [5:0] _GEN_38 = dType == 3'h3 ? 6'h1e : _GEN_13; // @[decode.scala 114:30 decode.scala 117:25]
  wire [63:0] _GEN_39 = dType == 3'h3 ? _dst_d_r_T : _GEN_31; // @[decode.scala 114:30 decode.scala 118:25]
  wire [63:0] _dst_d_r_T_6 = $signed(io_if2id_pc) + $signed(imm); // @[decode.scala 123:61]
  wire  _GEN_40 = dType == 3'h4 | _GEN_36; // @[decode.scala 120:30 decode.scala 121:25]
  wire  _GEN_41 = dType == 3'h4 | _GEN_37; // @[decode.scala 120:30 decode.scala 122:25]
  wire [63:0] _GEN_42 = dType == 3'h4 ? _dst_d_r_T_6 : _GEN_39; // @[decode.scala 120:30 decode.scala 123:25]
  wire [2:0] _GEN_43 = dType == 3'h4 ? io_if2id_inst[14:12] : ctrl_r_brType; // @[decode.scala 120:30 decode.scala 124:27 decode.scala 26:30]
  wire [1:0] _GEN_44 = dType == 3'h4 ? 2'h2 : _GEN_28; // @[decode.scala 120:30 decode.scala 125:25]
  wire [63:0] _GEN_45 = dType == 3'h5 ? _dst_d_r_T : _GEN_32; // @[decode.scala 127:30 decode.scala 128:25]
  wire [63:0] _GEN_46 = dType == 3'h5 ? io_if2id_pc : _GEN_30; // @[decode.scala 127:30 decode.scala 129:25]
  wire [63:0] _GEN_47 = dType == 3'h6 ? _dst_d_r_T_6 : _GEN_45; // @[decode.scala 131:30 decode.scala 132:25]
  wire [63:0] _GEN_48 = dType == 3'h6 ? _rs2_d_r_T_1 : _GEN_46; // @[decode.scala 131:30 decode.scala 133:25]
  wire [63:0] _GEN_49 = dType == 3'h6 ? 64'h0 : _GEN_42; // @[decode.scala 131:30 decode.scala 134:25]
  wire [1:0] _GEN_50 = dType == 3'h6 ? 2'h1 : _GEN_44; // @[decode.scala 131:30 decode.scala 135:24]
  wire  _excep_r_cause_T = io_idState_priv == 2'h3; // @[decode.scala 141:34]
  wire  _excep_r_cause_T_1 = io_idState_priv == 2'h1; // @[decode.scala 142:34]
  wire [3:0] _excep_r_cause_T_2 = _excep_r_cause_T_1 ? 4'h9 : 4'h8; // @[Mux.scala 47:69]
  wire [3:0] _excep_r_cause_T_3 = _excep_r_cause_T ? 4'hb : _excep_r_cause_T_2; // @[Mux.scala 47:69]
  wire [9:0] _rs2_r_T_4 = _excep_r_cause_T ? 10'h305 : 10'h105; // @[decode.scala 146:32]
  wire [63:0] _GEN_51 = 32'h73 == io_if2id_inst ? io_if2id_pc : _GEN_8; // @[decode.scala 137:38 decode.scala 138:25]
  wire  _GEN_52 = 32'h73 == io_if2id_inst | _GEN_5; // @[decode.scala 137:38 decode.scala 139:25]
  wire [63:0] _GEN_53 = 32'h73 == io_if2id_inst ? {{60'd0}, _excep_r_cause_T_3} : _GEN_6; // @[decode.scala 137:38 decode.scala 140:27]
  wire [63:0] _GEN_54 = 32'h73 == io_if2id_inst ? 64'h0 : _GEN_7; // @[decode.scala 137:38 decode.scala 144:27]
  wire [1:0] _GEN_55 = 32'h73 == io_if2id_inst ? 2'h3 : _GEN_50; // @[decode.scala 137:38 decode.scala 145:25]
  wire [11:0] _GEN_56 = 32'h73 == io_if2id_inst ? {{2'd0}, _rs2_r_T_4} : _rs2_r_T_2; // @[decode.scala 137:38 decode.scala 146:25 decode.scala 76:25]
  wire  _GEN_57 = 32'h73 == io_if2id_inst | _GEN_34; // @[decode.scala 137:38 decode.scala 43:17]
  wire  _GEN_58 = 32'h73 == io_if2id_inst | _GEN_35; // @[decode.scala 137:38 decode.scala 43:57]
  wire [63:0] _GEN_59 = 32'h10200073 == io_if2id_inst ? io_if2id_pc : _GEN_51; // @[decode.scala 149:37 decode.scala 150:25]
  wire  _GEN_60 = 32'h10200073 == io_if2id_inst | _GEN_52; // @[decode.scala 149:37 decode.scala 151:25]
  wire [1:0] _GEN_61 = 32'h10200073 == io_if2id_inst ? 2'h2 : 2'h0; // @[decode.scala 149:37 decode.scala 152:27]
  wire [63:0] _GEN_62 = 32'h10200073 == io_if2id_inst ? 64'h0 : _GEN_53; // @[decode.scala 149:37 decode.scala 153:27]
  wire [63:0] _GEN_63 = 32'h10200073 == io_if2id_inst ? 64'h0 : _GEN_54; // @[decode.scala 149:37 decode.scala 154:27]
  wire [1:0] _GEN_64 = 32'h10200073 == io_if2id_inst ? 2'h3 : _GEN_55; // @[decode.scala 149:37 decode.scala 155:25]
  wire [11:0] _GEN_65 = 32'h10200073 == io_if2id_inst ? 12'h141 : _GEN_56; // @[decode.scala 149:37 decode.scala 156:25]
  wire  _GEN_66 = 32'h10200073 == io_if2id_inst | _GEN_57; // @[decode.scala 149:37 decode.scala 43:17]
  wire  _GEN_67 = 32'h10200073 == io_if2id_inst | _GEN_58; // @[decode.scala 149:37 decode.scala 43:57]
  wire [63:0] _GEN_68 = 32'h30200073 == io_if2id_inst ? io_if2id_pc : _GEN_59; // @[decode.scala 159:37 decode.scala 160:25]
  wire  _GEN_69 = 32'h30200073 == io_if2id_inst | _GEN_60; // @[decode.scala 159:37 decode.scala 161:25]
  wire [1:0] _GEN_70 = 32'h30200073 == io_if2id_inst ? 2'h3 : _GEN_61; // @[decode.scala 159:37 decode.scala 162:27]
  wire [63:0] _GEN_71 = 32'h30200073 == io_if2id_inst ? 64'h0 : _GEN_62; // @[decode.scala 159:37 decode.scala 163:27]
  wire [63:0] _GEN_72 = 32'h30200073 == io_if2id_inst ? 64'h0 : _GEN_63; // @[decode.scala 159:37 decode.scala 164:27]
  wire [1:0] _GEN_73 = 32'h30200073 == io_if2id_inst ? 2'h3 : _GEN_64; // @[decode.scala 159:37 decode.scala 165:25]
  wire  _GEN_75 = 32'h30200073 == io_if2id_inst | _GEN_66; // @[decode.scala 159:37 decode.scala 43:17]
  wire  _GEN_76 = 32'h30200073 == io_if2id_inst | _GEN_67; // @[decode.scala 159:37 decode.scala 43:57]
  wire [1:0] _GEN_77 = _instType_T_183 ? 2'h1 : 2'h0; // @[decode.scala 169:40 decode.scala 170:23 decode.scala 80:25]
  wire  _GEN_78 = _instType_T_183 | _GEN_75; // @[decode.scala 169:40 decode.scala 43:17]
  wire  _GEN_79 = _instType_T_183 | _GEN_76; // @[decode.scala 169:40 decode.scala 43:57]
  wire [1:0] _GEN_80 = _instType_T_185 ? 2'h2 : _GEN_77; // @[decode.scala 173:43 decode.scala 174:23]
  wire  _GEN_81 = _instType_T_185 | _GEN_78; // @[decode.scala 173:43 decode.scala 43:17]
  wire  _GEN_82 = _instType_T_185 | _GEN_79; // @[decode.scala 173:43 decode.scala 43:57]
  wire  _GEN_105 = hs_in & ~is_compress & ~io_if2id_excep_en & _GEN_81; // @[decode.scala 65:54 decode.scala 19:33]
  wire [63:0] _GEN_106 = hs_in & ~is_compress & ~io_if2id_excep_en ? _GEN_48 : rs2_d_r; // @[decode.scala 65:54 decode.scala 32:30]
  wire [63:0] _GEN_107 = hs_in & ~is_compress & ~io_if2id_excep_en ? _GEN_49 : dst_d_r; // @[decode.scala 65:54 decode.scala 34:30]
  wire [63:0] _GEN_108 = hs_in & ~is_compress & ~io_if2id_excep_en ? _GEN_47 : rs1_d_r; // @[decode.scala 65:54 decode.scala 29:30]
  wire [2:0] _GEN_109 = hs_in & ~is_compress & ~io_if2id_excep_en ? _GEN_43 : ctrl_r_brType; // @[decode.scala 65:54 decode.scala 26:30]
  wire  _T_28 = 4'h1 == instType_c_1; // @[Conditional.scala 37:30]
  wire [3:0] imm_c_hi_hi_lo = io_if2id_inst[10:7]; // @[decode.scala 185:51]
  wire [1:0] imm_c_hi_lo = io_if2id_inst[12:11]; // @[decode.scala 185:65]
  wire  imm_c_lo_hi_hi = io_if2id_inst[5]; // @[decode.scala 185:80]
  wire  imm_c_lo_hi_lo = io_if2id_inst[6]; // @[decode.scala 185:91]
  wire [63:0] _imm_c_T_1 = {54'h0,imm_c_hi_hi_lo,imm_c_hi_lo,imm_c_lo_hi_hi,imm_c_lo_hi_lo,2'h0}; // @[decode.scala 185:106]
  wire  _T_29 = 4'h2 == instType_c_1; // @[Conditional.scala 37:30]
  wire [2:0] imm_c_hi_lo_1 = io_if2id_inst[12:10]; // @[decode.scala 186:62]
  wire [63:0] _imm_c_T_3 = {57'h0,imm_c_lo_hi_hi,imm_c_hi_lo_1,imm_c_lo_hi_lo,2'h0}; // @[decode.scala 186:92]
  wire  _T_30 = 4'h3 == instType_c_1; // @[Conditional.scala 37:30]
  wire [1:0] imm_c_hi_lo_2 = io_if2id_inst[6:5]; // @[decode.scala 187:51]
  wire [63:0] _imm_c_T_5 = {56'h0,imm_c_hi_lo_2,imm_c_hi_lo_1,3'h0}; // @[decode.scala 187:83]
  wire  _T_31 = 4'h4 == instType_c_1; // @[Conditional.scala 37:30]
  wire  imm_c_hi_lo_3 = io_if2id_inst[12]; // @[decode.scala 188:51]
  wire [4:0] imm_c_lo_3 = io_if2id_inst[6:2]; // @[decode.scala 188:63]
  wire [63:0] _imm_c_T_7 = {58'h0,imm_c_hi_lo_3,imm_c_lo_3}; // @[decode.scala 188:70]
  wire  _T_32 = 4'h5 == instType_c_1; // @[Conditional.scala 37:30]
  wire [5:0] _imm_c_T_9 = {imm_c_hi_lo_3,imm_c_lo_3}; // @[decode.scala 189:59]
  wire  _T_33 = 4'h6 == instType_c_1; // @[Conditional.scala 37:30]
  wire [1:0] imm_c_hi_hi_lo_2 = io_if2id_inst[3:2]; // @[decode.scala 190:51]
  wire [2:0] imm_c_lo_hi_3 = io_if2id_inst[6:4]; // @[decode.scala 190:76]
  wire [63:0] _imm_c_T_11 = {56'h0,imm_c_hi_hi_lo_2,imm_c_hi_lo_3,imm_c_lo_hi_3,2'h0}; // @[decode.scala 190:93]
  wire  _T_34 = 4'h7 == instType_c_1; // @[Conditional.scala 37:30]
  wire [2:0] imm_c_hi_hi_lo_3 = io_if2id_inst[4:2]; // @[decode.scala 191:51]
  wire [63:0] _imm_c_T_13 = {55'h0,imm_c_hi_hi_lo_3,imm_c_hi_lo_3,imm_c_hi_lo_2,3'h0}; // @[decode.scala 191:93]
  wire  _T_35 = 4'h8 == instType_c_1; // @[Conditional.scala 37:30]
  wire [1:0] imm_c_hi_hi_lo_4 = io_if2id_inst[4:3]; // @[decode.scala 192:52]
  wire  imm_c_lo_hi_hi_1 = io_if2id_inst[2]; // @[decode.scala 192:76]
  wire [9:0] _imm_c_T_15 = {imm_c_hi_lo_3,imm_c_hi_hi_lo_4,imm_c_lo_hi_hi,imm_c_lo_hi_hi_1,imm_c_lo_hi_lo,4'h0}; // @[decode.scala 192:102]
  wire  _T_36 = 4'h9 == instType_c_1; // @[Conditional.scala 37:30]
  wire [17:0] _imm_c_T_17 = {imm_c_hi_lo_3,imm_c_lo_3,12'h0}; // @[decode.scala 193:70]
  wire  _T_37 = 4'ha == instType_c_1; // @[Conditional.scala 37:30]
  wire  imm_c_hi_hi_hi_lo = io_if2id_inst[8]; // @[decode.scala 194:52]
  wire [1:0] imm_c_hi_hi_lo_5 = io_if2id_inst[10:9]; // @[decode.scala 194:63]
  wire  imm_c_hi_lo_lo = io_if2id_inst[7]; // @[decode.scala 194:88]
  wire  imm_c_lo_hi_lo_2 = io_if2id_inst[11]; // @[decode.scala 194:110]
  wire [2:0] imm_c_lo_lo_hi = io_if2id_inst[5:3]; // @[decode.scala 194:122]
  wire [11:0] _imm_c_T_19 = {imm_c_hi_lo_3,imm_c_hi_hi_hi_lo,imm_c_hi_hi_lo_5,imm_c_lo_hi_lo,imm_c_hi_lo_lo,
    imm_c_lo_hi_hi_1,imm_c_lo_hi_lo_2,imm_c_lo_lo_hi,1'h0}; // @[decode.scala 194:139]
  wire  _T_38 = 4'hb == instType_c_1; // @[Conditional.scala 37:30]
  wire [1:0] imm_c_lo_hi_hi_3 = io_if2id_inst[11:10]; // @[decode.scala 195:76]
  wire [8:0] _imm_c_T_21 = {imm_c_hi_lo_3,imm_c_hi_lo_2,imm_c_lo_hi_hi_1,imm_c_lo_hi_hi_3,imm_c_hi_hi_lo_4,1'h0}; // @[decode.scala 195:108]
  wire  _T_39 = 4'hc == instType_c_1; // @[Conditional.scala 37:30]
  wire [1:0] imm_c_hi_lo_10 = io_if2id_inst[8:7]; // @[decode.scala 196:51]
  wire [3:0] imm_c_lo_hi_8 = io_if2id_inst[12:9]; // @[decode.scala 196:64]
  wire [63:0] _imm_c_T_23 = {56'h0,imm_c_hi_lo_10,imm_c_lo_hi_8,2'h0}; // @[decode.scala 196:82]
  wire  _T_40 = 4'hd == instType_c_1; // @[Conditional.scala 37:30]
  wire [2:0] imm_c_hi_lo_11 = io_if2id_inst[9:7]; // @[decode.scala 197:51]
  wire [63:0] _imm_c_T_25 = {55'h0,imm_c_hi_lo_11,imm_c_hi_lo_1,3'h0}; // @[decode.scala 197:83]
  wire [63:0] _GEN_110 = _T_40 ? $signed(_imm_c_T_25) : $signed(64'sh0); // @[Conditional.scala 39:67 decode.scala 197:27 decode.scala 182:11]
  wire [63:0] _GEN_111 = _T_39 ? $signed(_imm_c_T_23) : $signed(_GEN_110); // @[Conditional.scala 39:67 decode.scala 196:27]
  wire [63:0] _GEN_112 = _T_38 ? $signed({{55{_imm_c_T_21[8]}},_imm_c_T_21}) : $signed(_GEN_111); // @[Conditional.scala 39:67 decode.scala 195:27]
  wire [63:0] _GEN_113 = _T_37 ? $signed({{52{_imm_c_T_19[11]}},_imm_c_T_19}) : $signed(_GEN_112); // @[Conditional.scala 39:67 decode.scala 194:27]
  wire [63:0] _GEN_114 = _T_36 ? $signed({{46{_imm_c_T_17[17]}},_imm_c_T_17}) : $signed(_GEN_113); // @[Conditional.scala 39:67 decode.scala 193:27]
  wire [63:0] _GEN_115 = _T_35 ? $signed({{54{_imm_c_T_15[9]}},_imm_c_T_15}) : $signed(_GEN_114); // @[Conditional.scala 39:67 decode.scala 192:27]
  wire [63:0] _GEN_116 = _T_34 ? $signed(_imm_c_T_13) : $signed(_GEN_115); // @[Conditional.scala 39:67 decode.scala 191:27]
  wire [63:0] _GEN_117 = _T_33 ? $signed(_imm_c_T_11) : $signed(_GEN_116); // @[Conditional.scala 39:67 decode.scala 190:27]
  wire [63:0] _GEN_118 = _T_32 ? $signed({{58{_imm_c_T_9[5]}},_imm_c_T_9}) : $signed(_GEN_117); // @[Conditional.scala 39:67 decode.scala 189:27]
  wire [63:0] _GEN_119 = _T_31 ? $signed(_imm_c_T_7) : $signed(_GEN_118); // @[Conditional.scala 39:67 decode.scala 188:27]
  wire [63:0] _GEN_120 = _T_30 ? $signed(_imm_c_T_5) : $signed(_GEN_119); // @[Conditional.scala 39:67 decode.scala 187:27]
  wire [63:0] _GEN_121 = _T_29 ? $signed(_imm_c_T_3) : $signed(_GEN_120); // @[Conditional.scala 39:67 decode.scala 186:27]
  wire [63:0] imm_c = _T_28 ? $signed(_imm_c_T_1) : $signed(_GEN_121); // @[Conditional.scala 40:58 decode.scala 185:27]
  wire [30:0] _inst_r_T = {15'h0,io_if2id_inst[15:0]}; // @[Cat.scala 30:58]
  wire  _GEN_123 = instType_c_0 == 4'h0 & _T_7 | io_if2id_excep_en; // @[decode.scala 218:58 decode.scala 219:29 decode.scala 202:25]
  wire  _GEN_128 = instType_c_0 == 4'h0 & _T_7 | _GEN_105; // @[decode.scala 218:58 decode.scala 43:17]
  wire  _GEN_129 = instType_c_0 == 4'h0 & _T_7 | io_if2id_recov; // @[decode.scala 218:58 decode.scala 43:57 decode.scala 217:25]
  wire  _T_47 = instType_c_0 == 4'h1; // @[decode.scala 226:22]
  wire [1:0] _GEN_130 = _instType_c_T_52 ? 2'h1 : 2'h0; // @[decode.scala 229:34 decode.scala 230:29 decode.scala 213:25]
  wire [63:0] _GEN_131 = _instType_c_T_52 ? 64'h0 : _GEN_107; // @[decode.scala 229:34 decode.scala 231:29]
  wire [63:0] _rs2_d_r_T_6 = io_if2id_pc + 64'h2; // @[decode.scala 236:44]
  wire [1:0] _GEN_132 = _instType_c_T_56 ? 2'h1 : _GEN_130; // @[decode.scala 233:36 decode.scala 234:29]
  wire  _GEN_133 = _instType_c_T_56 ? 1'h0 : 1'h1; // @[decode.scala 233:36 decode.scala 235:29 decode.scala 228:20]
  wire [63:0] _GEN_134 = _instType_c_T_56 ? _rs2_d_r_T_6 : _GEN_106; // @[decode.scala 233:36 decode.scala 236:29]
  wire [63:0] _GEN_135 = _instType_c_T_56 ? 64'h0 : _GEN_131; // @[decode.scala 233:36 decode.scala 237:29]
  wire [4:0] _GEN_136 = _instType_c_T_56 ? 5'h1 : io_if2id_inst[11:7]; // @[decode.scala 233:36 decode.scala 238:29 decode.scala 212:25]
  wire  _GEN_138 = instType_c_0 == 4'h1 & _GEN_133; // @[decode.scala 226:29 decode.scala 211:25]
  wire [1:0] _GEN_139 = instType_c_0 == 4'h1 ? _GEN_132 : 2'h0; // @[decode.scala 226:29 decode.scala 213:25]
  wire [63:0] _GEN_140 = instType_c_0 == 4'h1 ? _GEN_135 : _GEN_107; // @[decode.scala 226:29]
  wire [63:0] _GEN_141 = instType_c_0 == 4'h1 ? _GEN_134 : _GEN_106; // @[decode.scala 226:29]
  wire [4:0] _GEN_142 = instType_c_0 == 4'h1 ? _GEN_136 : io_if2id_inst[11:7]; // @[decode.scala 226:29 decode.scala 212:25]
  wire [63:0] _rs2_d_r_T_7 = _T_28 ? $signed(_imm_c_T_1) : $signed(_GEN_121); // @[decode.scala 243:30]
  wire [4:0] _GEN_143 = _instType_c_T_48 | _instType_c_T_50 ? 5'h2 : io_if2id_inst[11:7]; // @[decode.scala 244:57 decode.scala 245:23 decode.scala 208:25]
  wire  _GEN_144 = instType_c_0 == 4'h2 | _T_47; // @[decode.scala 241:29 decode.scala 242:21]
  wire [63:0] _GEN_145 = instType_c_0 == 4'h2 ? _rs2_d_r_T_7 : _GEN_141; // @[decode.scala 241:29 decode.scala 243:21]
  wire [4:0] _GEN_146 = instType_c_0 == 4'h2 ? _GEN_143 : io_if2id_inst[11:7]; // @[decode.scala 241:29 decode.scala 208:25]
  wire  _GEN_147 = instType_c_0 == 4'h3 | _GEN_144; // @[decode.scala 248:30 decode.scala 249:21]
  wire [4:0] _GEN_148 = instType_c_0 == 4'h3 ? 5'h2 : _GEN_146; // @[decode.scala 248:30 decode.scala 250:21]
  wire  _GEN_149 = instType_c_0 == 4'h3 | _GEN_138; // @[decode.scala 248:30 decode.scala 251:21]
  wire [4:0] _GEN_150 = instType_c_0 == 4'h3 ? imm_c_lo_3 : imm_c_lo_3; // @[decode.scala 248:30 decode.scala 252:21 decode.scala 210:25]
  wire [63:0] _GEN_151 = instType_c_0 == 4'h3 ? _rs2_d_r_T_7 : _GEN_140; // @[decode.scala 248:30 decode.scala 253:21]
  wire [5:0] _GEN_152 = instType_c_0 == 4'h3 ? 6'h1e : 6'h1b; // @[decode.scala 248:30 decode.scala 254:21 decode.scala 216:25]
  wire [3:0] _dst_r_T_3 = {1'h1,imm_c_hi_hi_lo_3}; // @[Cat.scala 30:58]
  wire  _GEN_153 = instType_c_0 == 4'h4 | _GEN_147; // @[decode.scala 256:30 decode.scala 257:21]
  wire [4:0] _GEN_154 = instType_c_0 == 4'h4 ? 5'h2 : _GEN_148; // @[decode.scala 256:30 decode.scala 258:21]
  wire [63:0] _GEN_155 = instType_c_0 == 4'h4 ? _rs2_d_r_T_7 : _GEN_145; // @[decode.scala 256:30 decode.scala 259:21]
  wire [4:0] _GEN_156 = instType_c_0 == 4'h4 ? {{1'd0}, _dst_r_T_3} : _GEN_142; // @[decode.scala 256:30 decode.scala 260:21]
  wire [3:0] _rs1_r_T_3 = {1'h1,imm_c_hi_lo_11}; // @[Cat.scala 30:58]
  wire  _GEN_157 = instType_c_0 == 4'h5 | _GEN_153; // @[decode.scala 262:29 decode.scala 263:21]
  wire [4:0] _GEN_158 = instType_c_0 == 4'h5 ? {{1'd0}, _rs1_r_T_3} : _GEN_154; // @[decode.scala 262:29 decode.scala 264:21]
  wire [4:0] _GEN_160 = instType_c_0 == 4'h5 ? {{1'd0}, _dst_r_T_3} : _GEN_156; // @[decode.scala 262:29 decode.scala 266:21]
  wire [5:0] _GEN_161 = io_if2id_inst[1:0] == 2'h0 ? 6'h1e : _GEN_152; // @[decode.scala 275:38 decode.scala 276:25]
  wire  _GEN_162 = instType_c_0 == 4'h6 | _GEN_157; // @[decode.scala 268:29 decode.scala 269:21]
  wire  _GEN_164 = instType_c_0 == 4'h6 | _GEN_149; // @[decode.scala 268:29 decode.scala 271:21]
  wire [4:0] _GEN_165 = instType_c_0 == 4'h6 ? {{1'd0}, _dst_r_T_3} : _GEN_150; // @[decode.scala 268:29 decode.scala 272:21]
  wire [63:0] _GEN_166 = instType_c_0 == 4'h6 ? _rs2_d_r_T_7 : _GEN_151; // @[decode.scala 268:29 decode.scala 273:21]
  wire [63:0] _dst_d_r_T_13 = $signed(io_if2id_pc) + $signed(imm_c); // @[decode.scala 283:53]
  wire [2:0] _GEN_169 = _instType_c_T_42 ? 3'h0 : _GEN_109; // @[decode.scala 285:36 decode.scala 286:31]
  wire [63:0] _GEN_170 = _instType_c_T_42 ? 64'h0 : _rs2_d_r_T_7; // @[decode.scala 285:36 decode.scala 287:29 decode.scala 282:21]
  wire [1:0] _GEN_171 = _instType_c_T_42 ? 2'h2 : _GEN_139; // @[decode.scala 285:36 decode.scala 288:29]
  wire [2:0] _GEN_172 = _instType_c_T_44 ? 3'h1 : _GEN_169; // @[decode.scala 290:36 decode.scala 291:31]
  wire [1:0] _GEN_174 = _instType_c_T_44 ? 2'h2 : _GEN_171; // @[decode.scala 290:36 decode.scala 293:29]
  wire  _GEN_175 = instType_c_0 == 4'h7 | _GEN_162; // @[decode.scala 279:29 decode.scala 280:21]
  wire [1:0] _GEN_181 = instType_c_0 == 4'h7 ? _GEN_174 : _GEN_139; // @[decode.scala 279:29]
  wire  _GEN_233 = valid_r & ~hs_out ? 1'h0 : io_if2id_valid; // @[decode.scala 318:33 decode.scala 316:20]
  wire  _GEN_235 = hs_out ? 1'h0 : valid_r; // @[decode.scala 326:26 decode.scala 327:20 decode.scala 40:30]
  wire  _GEN_236 = hs_in | _GEN_235; // @[decode.scala 324:19 decode.scala 325:20]
  wire  _GEN_237 = _io_if2id_stall_T & _GEN_236; // @[decode.scala 323:25 decode.scala 331:17]
  assign io_if2id_drop = drop_r | io_id2df_drop; // @[decode.scala 20:30]
  assign io_if2id_stall = stall_r & ~io_id2df_drop | io_id2df_stall; // @[decode.scala 22:52]
  assign io_if2id_ready = ~drop_in & _GEN_233; // @[decode.scala 317:19 decode.scala 316:20]
  assign io_id2df_inst = inst_r; // @[decode.scala 333:25]
  assign io_id2df_pc = pc_r; // @[decode.scala 334:25]
  assign io_id2df_excep_cause = excep_r_cause; // @[decode.scala 335:25]
  assign io_id2df_excep_tval = excep_r_tval; // @[decode.scala 335:25]
  assign io_id2df_excep_en = excep_r_en; // @[decode.scala 335:25]
  assign io_id2df_excep_pc = excep_r_pc; // @[decode.scala 335:25]
  assign io_id2df_excep_etype = excep_r_etype; // @[decode.scala 335:25]
  assign io_id2df_ctrl_aluOp = ctrl_r_aluOp; // @[decode.scala 336:25]
  assign io_id2df_ctrl_aluWidth = ctrl_r_aluWidth; // @[decode.scala 336:25]
  assign io_id2df_ctrl_dcMode = ctrl_r_dcMode; // @[decode.scala 336:25]
  assign io_id2df_ctrl_writeRegEn = ctrl_r_writeRegEn; // @[decode.scala 336:25]
  assign io_id2df_ctrl_writeCSREn = ctrl_r_writeCSREn; // @[decode.scala 336:25]
  assign io_id2df_ctrl_brType = ctrl_r_brType; // @[decode.scala 336:25]
  assign io_id2df_rs1 = rs1_r; // @[decode.scala 337:25]
  assign io_id2df_rrs1 = rrs1_r; // @[decode.scala 338:25]
  assign io_id2df_rs1_d = rs1_d_r; // @[decode.scala 339:25]
  assign io_id2df_rs2 = rs2_r; // @[decode.scala 340:25]
  assign io_id2df_rrs2 = rrs2_r; // @[decode.scala 341:25]
  assign io_id2df_rs2_d = rs2_d_r; // @[decode.scala 342:25]
  assign io_id2df_dst = dst_r; // @[decode.scala 343:25]
  assign io_id2df_dst_d = dst_d_r; // @[decode.scala 344:25]
  assign io_id2df_jmp_type = jmp_type_r; // @[decode.scala 345:25]
  assign io_id2df_special = special_r; // @[decode.scala 346:25]
  assign io_id2df_swap = swap_r; // @[decode.scala 347:25]
  assign io_id2df_indi = indi_r; // @[decode.scala 348:25]
  assign io_id2df_recov = recov_r; // @[decode.scala 349:25]
  assign io_id2df_valid = valid_r; // @[decode.scala 350:25]
  always @(posedge clock) begin
    if (reset) begin // @[decode.scala 17:30]
      drop_r <= 1'h0; // @[decode.scala 17:30]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      drop_r <= _GEN_128;
    end else begin
      drop_r <= _GEN_105;
    end
    if (reset) begin // @[decode.scala 18:30]
      stall_r <= 1'h0; // @[decode.scala 18:30]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      stall_r <= _GEN_128;
    end else begin
      stall_r <= _GEN_105;
    end
    if (reset) begin // @[decode.scala 23:30]
      inst_r <= 32'h0; // @[decode.scala 23:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      inst_r <= io_if2id_inst; // @[decode.scala 303:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      inst_r <= {{1'd0}, _inst_r_T}; // @[decode.scala 200:17]
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      inst_r <= io_if2id_inst; // @[decode.scala 66:25]
    end
    if (reset) begin // @[decode.scala 24:30]
      pc_r <= 64'h0; // @[decode.scala 24:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      pc_r <= io_if2id_pc; // @[decode.scala 304:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      pc_r <= io_if2id_pc; // @[decode.scala 201:17]
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      pc_r <= io_if2id_pc; // @[decode.scala 67:25]
    end
    if (reset) begin // @[decode.scala 25:30]
      excep_r_cause <= 64'h0; // @[decode.scala 25:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      excep_r_cause <= io_if2id_excep_cause; // @[decode.scala 305:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      if (instType_c_0 == 4'h0 & _T_7) begin // @[decode.scala 218:58]
        excep_r_cause <= 64'h2; // @[decode.scala 220:29]
      end else begin
        excep_r_cause <= io_if2id_excep_cause; // @[decode.scala 202:25]
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      excep_r_cause <= _GEN_71;
    end
    if (reset) begin // @[decode.scala 25:30]
      excep_r_tval <= 64'h0; // @[decode.scala 25:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      excep_r_tval <= io_if2id_excep_tval; // @[decode.scala 305:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      if (instType_c_0 == 4'h0 & _T_7) begin // @[decode.scala 218:58]
        excep_r_tval <= {{33'd0}, _inst_r_T}; // @[decode.scala 221:29]
      end else begin
        excep_r_tval <= io_if2id_excep_tval; // @[decode.scala 202:25]
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      excep_r_tval <= _GEN_72;
    end
    if (reset) begin // @[decode.scala 25:30]
      excep_r_en <= 1'h0; // @[decode.scala 25:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      excep_r_en <= io_if2id_excep_en; // @[decode.scala 305:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      excep_r_en <= _GEN_123;
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      excep_r_en <= _GEN_69;
    end
    if (reset) begin // @[decode.scala 25:30]
      excep_r_pc <= 64'h0; // @[decode.scala 25:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      excep_r_pc <= io_if2id_excep_pc; // @[decode.scala 305:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      if (instType_c_0 == 4'h0 & _T_7) begin // @[decode.scala 218:58]
        excep_r_pc <= io_if2id_pc; // @[decode.scala 222:29]
      end else begin
        excep_r_pc <= io_if2id_excep_pc; // @[decode.scala 202:25]
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      excep_r_pc <= _GEN_68;
    end
    if (reset) begin // @[decode.scala 25:30]
      excep_r_etype <= 2'h0; // @[decode.scala 25:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      excep_r_etype <= 2'h0; // @[decode.scala 305:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      excep_r_etype <= 2'h0;
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      excep_r_etype <= _GEN_70;
    end
    if (reset) begin // @[decode.scala 26:30]
      ctrl_r_aluOp <= 5'h0; // @[decode.scala 26:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      ctrl_r_aluOp <= 5'h0; // @[decode.scala 306:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      if (_instType_c_T_2) begin // @[Lookup.scala 33:37]
        ctrl_r_aluOp <= 5'h3;
      end else begin
        ctrl_r_aluOp <= _instType_c_T_152;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      ctrl_r_aluOp <= instType_1; // @[decode.scala 69:27]
    end
    if (reset) begin // @[decode.scala 26:30]
      ctrl_r_aluWidth <= 1'h0; // @[decode.scala 26:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      ctrl_r_aluWidth <= 1'h0; // @[decode.scala 306:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      if (_instType_c_T_2) begin // @[Lookup.scala 33:37]
        ctrl_r_aluWidth <= 1'h0;
      end else begin
        ctrl_r_aluWidth <= _instType_c_T_182;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      ctrl_r_aluWidth <= instType_2; // @[decode.scala 70:27]
    end
    if (reset) begin // @[decode.scala 26:30]
      ctrl_r_dcMode <= 5'h0; // @[decode.scala 26:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      ctrl_r_dcMode <= 5'h0; // @[decode.scala 306:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      if (_instType_c_T_2) begin // @[Lookup.scala 33:37]
        ctrl_r_dcMode <= 5'h0;
      end else begin
        ctrl_r_dcMode <= _instType_c_T_212;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      ctrl_r_dcMode <= instType_3; // @[decode.scala 71:27]
    end
    if (reset) begin // @[decode.scala 26:30]
      ctrl_r_writeRegEn <= 1'h0; // @[decode.scala 26:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      ctrl_r_writeRegEn <= 1'h0; // @[decode.scala 306:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      ctrl_r_writeRegEn <= instType_c_5; // @[decode.scala 206:27]
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      ctrl_r_writeRegEn <= instType_4; // @[decode.scala 72:27]
    end
    if (reset) begin // @[decode.scala 26:30]
      ctrl_r_writeCSREn <= 1'h0; // @[decode.scala 26:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      ctrl_r_writeCSREn <= 1'h0; // @[decode.scala 306:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      ctrl_r_writeCSREn <= 1'h0; // @[decode.scala 207:27]
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      ctrl_r_writeCSREn <= instType_6; // @[decode.scala 73:27]
    end
    if (reset) begin // @[decode.scala 26:30]
      ctrl_r_brType <= 3'h0; // @[decode.scala 26:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      ctrl_r_brType <= 3'h0; // @[decode.scala 306:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      if (instType_c_0 == 4'h7) begin // @[decode.scala 279:29]
        ctrl_r_brType <= _GEN_172;
      end else begin
        ctrl_r_brType <= _GEN_109;
      end
    end else begin
      ctrl_r_brType <= _GEN_109;
    end
    if (reset) begin // @[decode.scala 27:30]
      rs1_r <= 5'h0; // @[decode.scala 27:30]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      if (instType_c_0 == 4'h7) begin // @[decode.scala 279:29]
        rs1_r <= {{1'd0}, _rs1_r_T_3}; // @[decode.scala 281:21]
      end else if (instType_c_0 == 4'h6) begin // @[decode.scala 268:29]
        rs1_r <= {{1'd0}, _rs1_r_T_3}; // @[decode.scala 270:21]
      end else begin
        rs1_r <= _GEN_158;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      rs1_r <= io_if2id_inst[19:15]; // @[decode.scala 74:25]
    end
    if (reset) begin // @[decode.scala 28:30]
      rrs1_r <= 1'h0; // @[decode.scala 28:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      rrs1_r <= 1'h0; // @[decode.scala 307:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      rrs1_r <= _GEN_175;
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      rrs1_r <= _GEN_40;
    end
    if (reset) begin // @[decode.scala 29:30]
      rs1_d_r <= 64'h0; // @[decode.scala 29:30]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      if (instType_c_0 == 4'h8) begin // @[decode.scala 296:29]
        rs1_d_r <= io_if2id_pc; // @[decode.scala 297:21]
      end else begin
        rs1_d_r <= _GEN_108;
      end
    end else begin
      rs1_d_r <= _GEN_108;
    end
    if (reset) begin // @[decode.scala 30:30]
      rs2_r <= 12'h0; // @[decode.scala 30:30]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      rs2_r <= {{7'd0}, _GEN_165};
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      if (32'h30200073 == io_if2id_inst) begin // @[decode.scala 159:37]
        rs2_r <= 12'h341; // @[decode.scala 166:25]
      end else begin
        rs2_r <= _GEN_65;
      end
    end
    if (reset) begin // @[decode.scala 31:30]
      rrs2_r <= 1'h0; // @[decode.scala 31:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      rrs2_r <= 1'h0; // @[decode.scala 308:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      rrs2_r <= _GEN_164;
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      rrs2_r <= _GEN_41;
    end
    if (reset) begin // @[decode.scala 32:30]
      rs2_d_r <= 64'h0; // @[decode.scala 32:30]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      if (instType_c_0 == 4'h7) begin // @[decode.scala 279:29]
        if (_instType_c_T_44) begin // @[decode.scala 290:36]
          rs2_d_r <= 64'h0; // @[decode.scala 292:29]
        end else begin
          rs2_d_r <= _GEN_170;
        end
      end else if (instType_c_0 == 4'h5) begin // @[decode.scala 262:29]
        rs2_d_r <= _rs2_d_r_T_7; // @[decode.scala 265:21]
      end else begin
        rs2_d_r <= _GEN_155;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      if (dType == 3'h6) begin // @[decode.scala 131:30]
        rs2_d_r <= _rs2_d_r_T_1; // @[decode.scala 133:25]
      end else begin
        rs2_d_r <= _GEN_46;
      end
    end
    if (reset) begin // @[decode.scala 33:30]
      dst_r <= 5'h0; // @[decode.scala 33:30]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      if (instType_c_0 == 4'h7) begin // @[decode.scala 279:29]
        dst_r <= {{1'd0}, _rs1_r_T_3}; // @[decode.scala 284:21]
      end else if (instType_c_0 == 4'h6) begin // @[decode.scala 268:29]
        dst_r <= {{1'd0}, _rs1_r_T_3}; // @[decode.scala 274:21]
      end else begin
        dst_r <= _GEN_160;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      dst_r <= imm_lo; // @[decode.scala 78:25]
    end
    if (reset) begin // @[decode.scala 34:30]
      dst_d_r <= 64'h0; // @[decode.scala 34:30]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      if (instType_c_0 == 4'h8) begin // @[decode.scala 296:29]
        dst_d_r <= _rs2_d_r_T_7; // @[decode.scala 298:21]
      end else if (instType_c_0 == 4'h7) begin // @[decode.scala 279:29]
        dst_d_r <= _dst_d_r_T_13; // @[decode.scala 283:21]
      end else begin
        dst_d_r <= _GEN_166;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      if (dType == 3'h6) begin // @[decode.scala 131:30]
        dst_d_r <= 64'h0; // @[decode.scala 134:25]
      end else begin
        dst_d_r <= _GEN_42;
      end
    end
    if (reset) begin // @[decode.scala 35:30]
      jmp_type_r <= 2'h0; // @[decode.scala 35:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      jmp_type_r <= 2'h0; // @[decode.scala 309:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      if (instType_c_0 == 4'h8) begin // @[decode.scala 296:29]
        jmp_type_r <= 2'h1; // @[decode.scala 299:25]
      end else begin
        jmp_type_r <= _GEN_181;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      jmp_type_r <= _GEN_73;
    end
    if (reset) begin // @[decode.scala 36:30]
      special_r <= 2'h0; // @[decode.scala 36:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      special_r <= 2'h0; // @[decode.scala 310:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      special_r <= 2'h0; // @[decode.scala 214:25]
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      special_r <= _GEN_80;
    end
    if (reset) begin // @[decode.scala 37:30]
      swap_r <= 6'h0; // @[decode.scala 37:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      swap_r <= 6'h1b; // @[decode.scala 312:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      if (instType_c_0 == 4'h6) begin // @[decode.scala 268:29]
        swap_r <= _GEN_161;
      end else begin
        swap_r <= _GEN_152;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      swap_r <= _GEN_38;
    end
    if (reset) begin // @[decode.scala 38:30]
      indi_r <= 2'h0; // @[decode.scala 38:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      indi_r <= 2'h0; // @[decode.scala 311:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      indi_r <= 2'h0; // @[decode.scala 215:25]
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      indi_r <= _indi_r_T_8; // @[decode.scala 81:25]
    end
    if (reset) begin // @[decode.scala 39:30]
      recov_r <= 1'h0; // @[decode.scala 39:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[decode.scala 302:37]
      recov_r <= io_if2id_recov; // @[decode.scala 313:25]
    end else if (hs_in & is_compress & _T_7) begin // @[decode.scala 199:53]
      recov_r <= _GEN_129;
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[decode.scala 65:54]
      recov_r <= _GEN_82;
    end
    if (reset) begin // @[decode.scala 40:30]
      valid_r <= 1'h0; // @[decode.scala 40:30]
    end else begin
      valid_r <= _GEN_237;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  drop_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  stall_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  inst_r = _RAND_2[31:0];
  _RAND_3 = {2{`RANDOM}};
  pc_r = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  excep_r_cause = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  excep_r_tval = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  excep_r_en = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  excep_r_pc = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  excep_r_etype = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  ctrl_r_aluOp = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  ctrl_r_aluWidth = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ctrl_r_dcMode = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  ctrl_r_writeRegEn = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  ctrl_r_writeCSREn = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  ctrl_r_brType = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  rs1_r = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  rrs1_r = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  rs1_d_r = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  rs2_r = _RAND_18[11:0];
  _RAND_19 = {1{`RANDOM}};
  rrs2_r = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  rs2_d_r = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  dst_r = _RAND_21[4:0];
  _RAND_22 = {2{`RANDOM}};
  dst_d_r = _RAND_22[63:0];
  _RAND_23 = {1{`RANDOM}};
  jmp_type_r = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  special_r = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  swap_r = _RAND_25[5:0];
  _RAND_26 = {1{`RANDOM}};
  indi_r = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  recov_r = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_r = _RAND_28[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_Forwarding(
  input         clock,
  input         reset,
  input  [31:0] io_id2df_inst,
  input  [63:0] io_id2df_pc,
  input  [63:0] io_id2df_excep_cause,
  input  [63:0] io_id2df_excep_tval,
  input         io_id2df_excep_en,
  input  [63:0] io_id2df_excep_pc,
  input  [1:0]  io_id2df_excep_etype,
  input  [4:0]  io_id2df_ctrl_aluOp,
  input         io_id2df_ctrl_aluWidth,
  input  [4:0]  io_id2df_ctrl_dcMode,
  input         io_id2df_ctrl_writeRegEn,
  input         io_id2df_ctrl_writeCSREn,
  input  [2:0]  io_id2df_ctrl_brType,
  input  [4:0]  io_id2df_rs1,
  input         io_id2df_rrs1,
  input  [63:0] io_id2df_rs1_d,
  input  [11:0] io_id2df_rs2,
  input         io_id2df_rrs2,
  input  [63:0] io_id2df_rs2_d,
  input  [4:0]  io_id2df_dst,
  input  [63:0] io_id2df_dst_d,
  input  [1:0]  io_id2df_jmp_type,
  input  [1:0]  io_id2df_special,
  input  [5:0]  io_id2df_swap,
  input  [1:0]  io_id2df_indi,
  output        io_id2df_drop,
  output        io_id2df_stall,
  input         io_id2df_recov,
  input         io_id2df_valid,
  output        io_id2df_ready,
  output [31:0] io_df2rr_inst,
  output [63:0] io_df2rr_pc,
  output [63:0] io_df2rr_excep_cause,
  output [63:0] io_df2rr_excep_tval,
  output        io_df2rr_excep_en,
  output [63:0] io_df2rr_excep_pc,
  output [1:0]  io_df2rr_excep_etype,
  output [4:0]  io_df2rr_ctrl_aluOp,
  output        io_df2rr_ctrl_aluWidth,
  output [4:0]  io_df2rr_ctrl_dcMode,
  output        io_df2rr_ctrl_writeRegEn,
  output        io_df2rr_ctrl_writeCSREn,
  output [2:0]  io_df2rr_ctrl_brType,
  output [4:0]  io_df2rr_rs1,
  output        io_df2rr_rrs1,
  output [63:0] io_df2rr_rs1_d,
  output [11:0] io_df2rr_rs2,
  output        io_df2rr_rrs2,
  output [63:0] io_df2rr_rs2_d,
  output [4:0]  io_df2rr_dst,
  output [63:0] io_df2rr_dst_d,
  output [1:0]  io_df2rr_jmp_type,
  output [1:0]  io_df2rr_special,
  output [5:0]  io_df2rr_swap,
  output [1:0]  io_df2rr_indi,
  input         io_df2rr_drop,
  input         io_df2rr_stall,
  output        io_df2rr_recov,
  output        io_df2rr_valid,
  input         io_df2rr_ready,
  input  [4:0]  io_d_rr_id,
  input  [63:0] io_d_rr_data,
  input  [1:0]  io_d_rr_state,
  input  [4:0]  io_d_ex_id,
  input  [63:0] io_d_ex_data,
  input  [1:0]  io_d_ex_state,
  input  [4:0]  io_d_mem1_id,
  input  [63:0] io_d_mem1_data,
  input  [1:0]  io_d_mem1_state,
  input  [4:0]  io_d_mem2_id,
  input  [63:0] io_d_mem2_data,
  input  [1:0]  io_d_mem2_state,
  input  [4:0]  io_d_mem3_id,
  input  [63:0] io_d_mem3_data,
  input  [1:0]  io_d_mem3_state
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
`endif // RANDOMIZE_REG_INIT
  wire  _io_id2df_stall_T = ~io_df2rr_drop; // @[forwading.scala 23:36]
  reg [31:0] inst_r; // @[forwading.scala 24:30]
  reg [63:0] pc_r; // @[forwading.scala 25:30]
  reg [63:0] excep_r_cause; // @[forwading.scala 26:30]
  reg [63:0] excep_r_tval; // @[forwading.scala 26:30]
  reg  excep_r_en; // @[forwading.scala 26:30]
  reg [63:0] excep_r_pc; // @[forwading.scala 26:30]
  reg [1:0] excep_r_etype; // @[forwading.scala 26:30]
  reg [4:0] ctrl_r_aluOp; // @[forwading.scala 27:30]
  reg  ctrl_r_aluWidth; // @[forwading.scala 27:30]
  reg [4:0] ctrl_r_dcMode; // @[forwading.scala 27:30]
  reg  ctrl_r_writeRegEn; // @[forwading.scala 27:30]
  reg  ctrl_r_writeCSREn; // @[forwading.scala 27:30]
  reg [2:0] ctrl_r_brType; // @[forwading.scala 27:30]
  reg [4:0] rs1_r; // @[forwading.scala 28:30]
  reg  rrs1_r; // @[forwading.scala 29:30]
  reg [63:0] rs1_d_r; // @[forwading.scala 30:30]
  reg [11:0] rs2_r; // @[forwading.scala 31:30]
  reg  rrs2_r; // @[forwading.scala 32:30]
  reg [63:0] rs2_d_r; // @[forwading.scala 33:30]
  reg [4:0] dst_r; // @[forwading.scala 34:30]
  reg [63:0] dst_d_r; // @[forwading.scala 35:30]
  reg [1:0] jmp_type_r; // @[forwading.scala 36:30]
  reg [1:0] special_r; // @[forwading.scala 37:30]
  reg [1:0] indi_r; // @[forwading.scala 38:30]
  reg [5:0] swap_r; // @[forwading.scala 39:30]
  reg  recov_r; // @[forwading.scala 40:30]
  reg  valid_r; // @[forwading.scala 41:30]
  reg [4:0] pre_dst; // @[forwading.scala 43:30]
  reg  pre_wr; // @[forwading.scala 44:30]
  reg  state; // @[forwading.scala 47:24]
  wire  hs_in = io_id2df_ready & io_id2df_valid; // @[forwading.scala 48:34]
  wire  hs_out = io_df2rr_ready & io_df2rr_valid; // @[forwading.scala 49:34]
  wire [4:0] cur_rs1 = hs_in ? io_id2df_rs1 : rs1_r; // @[forwading.scala 59:26]
  wire  cur_rrs1 = hs_in ? io_id2df_rrs1 : rrs1_r; // @[forwading.scala 60:26]
  wire [11:0] cur_rs2 = hs_in ? io_id2df_rs2 : rs2_r; // @[forwading.scala 61:26]
  wire  cur_rrs2 = hs_in ? io_id2df_rrs2 : rrs2_r; // @[forwading.scala 62:26]
  wire  _T_1 = valid_r & pre_wr; // @[forwading.scala 67:28]
  wire  _T_5 = io_d_rr_state != 2'h0; // @[forwading.scala 69:63]
  wire  _T_7 = io_d_rr_state == 2'h1; // @[forwading.scala 70:32]
  wire [63:0] _GEN_0 = io_d_rr_state == 2'h1 ? io_d_rr_data : 64'h0; // @[forwading.scala 70:44 forwading.scala 71:26 forwading.scala 57:62]
  wire  _GEN_2 = io_d_rr_state == 2'h1 ? 1'h0 : 1'h1; // @[forwading.scala 70:44 forwading.scala 57:41 forwading.scala 74:26]
  wire  _T_9 = io_d_ex_state != 2'h0; // @[forwading.scala 76:63]
  wire  _T_11 = io_d_ex_state == 2'h1; // @[forwading.scala 77:32]
  wire [63:0] _GEN_3 = io_d_ex_state == 2'h1 ? io_d_ex_data : 64'h0; // @[forwading.scala 77:44 forwading.scala 78:26 forwading.scala 57:62]
  wire  _GEN_5 = io_d_ex_state == 2'h1 ? 1'h0 : 1'h1; // @[forwading.scala 77:44 forwading.scala 57:41 forwading.scala 81:26]
  wire  _T_13 = io_d_mem1_state != 2'h0; // @[forwading.scala 83:67]
  wire  _T_15 = io_d_mem1_state == 2'h1; // @[forwading.scala 84:34]
  wire [63:0] _GEN_6 = io_d_mem1_state == 2'h1 ? io_d_mem1_data : 64'h0; // @[forwading.scala 84:46 forwading.scala 85:26 forwading.scala 57:62]
  wire  _GEN_8 = io_d_mem1_state == 2'h1 ? 1'h0 : 1'h1; // @[forwading.scala 84:46 forwading.scala 57:41 forwading.scala 88:26]
  wire  _T_17 = io_d_mem2_state != 2'h0; // @[forwading.scala 90:67]
  wire  _T_19 = io_d_mem2_state == 2'h1; // @[forwading.scala 91:34]
  wire [63:0] _GEN_9 = io_d_mem2_state == 2'h1 ? io_d_mem2_data : 64'h0; // @[forwading.scala 91:46 forwading.scala 92:26 forwading.scala 57:62]
  wire  _GEN_11 = io_d_mem2_state == 2'h1 ? 1'h0 : 1'h1; // @[forwading.scala 91:46 forwading.scala 57:41 forwading.scala 95:26]
  wire  _T_21 = io_d_mem3_state != 2'h0; // @[forwading.scala 97:67]
  wire  _T_23 = io_d_mem3_state == 2'h1; // @[forwading.scala 98:34]
  wire [63:0] _GEN_12 = io_d_mem3_state == 2'h1 ? io_d_mem3_data : 64'h0; // @[forwading.scala 98:46 forwading.scala 99:26 forwading.scala 57:62]
  wire  _GEN_14 = io_d_mem3_state == 2'h1 ? 1'h0 : 1'h1; // @[forwading.scala 98:46 forwading.scala 57:41 forwading.scala 102:26]
  wire [63:0] _GEN_15 = cur_rs1 == io_d_mem3_id & io_d_mem3_state != 2'h0 ? _GEN_12 : 64'h0; // @[forwading.scala 97:82 forwading.scala 57:62]
  wire  _GEN_16 = cur_rs1 == io_d_mem3_id & io_d_mem3_state != 2'h0 & _T_23; // @[forwading.scala 97:82 forwading.scala 57:15]
  wire  _GEN_17 = cur_rs1 == io_d_mem3_id & io_d_mem3_state != 2'h0 & _GEN_14; // @[forwading.scala 97:82 forwading.scala 57:41]
  wire [63:0] _GEN_18 = cur_rs1 == io_d_mem2_id & io_d_mem2_state != 2'h0 ? _GEN_9 : _GEN_15; // @[forwading.scala 90:82]
  wire  _GEN_19 = cur_rs1 == io_d_mem2_id & io_d_mem2_state != 2'h0 ? _T_19 : _GEN_16; // @[forwading.scala 90:82]
  wire  _GEN_20 = cur_rs1 == io_d_mem2_id & io_d_mem2_state != 2'h0 ? _GEN_11 : _GEN_17; // @[forwading.scala 90:82]
  wire [63:0] _GEN_21 = cur_rs1 == io_d_mem1_id & io_d_mem1_state != 2'h0 ? _GEN_6 : _GEN_18; // @[forwading.scala 83:82]
  wire  _GEN_22 = cur_rs1 == io_d_mem1_id & io_d_mem1_state != 2'h0 ? _T_15 : _GEN_19; // @[forwading.scala 83:82]
  wire  _GEN_23 = cur_rs1 == io_d_mem1_id & io_d_mem1_state != 2'h0 ? _GEN_8 : _GEN_20; // @[forwading.scala 83:82]
  wire [63:0] _GEN_24 = cur_rs1 == io_d_ex_id & io_d_ex_state != 2'h0 ? _GEN_3 : _GEN_21; // @[forwading.scala 76:78]
  wire  _GEN_25 = cur_rs1 == io_d_ex_id & io_d_ex_state != 2'h0 ? _T_11 : _GEN_22; // @[forwading.scala 76:78]
  wire  _GEN_26 = cur_rs1 == io_d_ex_id & io_d_ex_state != 2'h0 ? _GEN_5 : _GEN_23; // @[forwading.scala 76:78]
  wire [63:0] _GEN_27 = cur_rs1 == io_d_rr_id & io_d_rr_state != 2'h0 ? _GEN_0 : _GEN_24; // @[forwading.scala 69:78]
  wire  _GEN_28 = cur_rs1 == io_d_rr_id & io_d_rr_state != 2'h0 ? _T_7 : _GEN_25; // @[forwading.scala 69:78]
  wire  _GEN_29 = cur_rs1 == io_d_rr_id & io_d_rr_state != 2'h0 ? _GEN_2 : _GEN_26; // @[forwading.scala 69:78]
  wire  _GEN_30 = valid_r & pre_wr & cur_rs1 == pre_dst | _GEN_29; // @[forwading.scala 67:59 forwading.scala 68:22]
  wire [63:0] _GEN_31 = valid_r & pre_wr & cur_rs1 == pre_dst ? 64'h0 : _GEN_27; // @[forwading.scala 67:59 forwading.scala 57:62]
  wire  _GEN_32 = valid_r & pre_wr & cur_rs1 == pre_dst ? 1'h0 : _GEN_28; // @[forwading.scala 67:59 forwading.scala 57:15]
  wire  _GEN_33 = cur_rs1 == 5'h0 ? 1'h0 : _GEN_30; // @[forwading.scala 65:30 forwading.scala 66:22]
  wire [63:0] _GEN_34 = cur_rs1 == 5'h0 ? 64'h0 : _GEN_31; // @[forwading.scala 65:30 forwading.scala 57:62]
  wire  _GEN_35 = cur_rs1 == 5'h0 ? 1'h0 : _GEN_32; // @[forwading.scala 65:30 forwading.scala 57:15]
  wire  rs1_wait = cur_rrs1 & _GEN_33; // @[forwading.scala 63:19 forwading.scala 57:41]
  wire  rs1_valid = cur_rrs1 & _GEN_35; // @[forwading.scala 63:19 forwading.scala 57:15]
  wire [11:0] _GEN_130 = {{7'd0}, pre_dst}; // @[forwading.scala 110:48]
  wire [11:0] _GEN_131 = {{7'd0}, io_d_rr_id}; // @[forwading.scala 112:29]
  wire [11:0] _GEN_132 = {{7'd0}, io_d_ex_id}; // @[forwading.scala 119:29]
  wire [11:0] _GEN_133 = {{7'd0}, io_d_mem1_id}; // @[forwading.scala 126:29]
  wire [11:0] _GEN_134 = {{7'd0}, io_d_mem2_id}; // @[forwading.scala 133:29]
  wire [11:0] _GEN_135 = {{7'd0}, io_d_mem3_id}; // @[forwading.scala 140:29]
  wire [63:0] _GEN_54 = cur_rs2 == _GEN_135 & _T_21 ? _GEN_12 : 64'h0; // @[forwading.scala 140:82 forwading.scala 58:62]
  wire  _GEN_55 = cur_rs2 == _GEN_135 & _T_21 & _T_23; // @[forwading.scala 140:82 forwading.scala 58:15]
  wire  _GEN_56 = cur_rs2 == _GEN_135 & _T_21 & _GEN_14; // @[forwading.scala 140:82 forwading.scala 58:41]
  wire [63:0] _GEN_57 = cur_rs2 == _GEN_134 & _T_17 ? _GEN_9 : _GEN_54; // @[forwading.scala 133:82]
  wire  _GEN_58 = cur_rs2 == _GEN_134 & _T_17 ? _T_19 : _GEN_55; // @[forwading.scala 133:82]
  wire  _GEN_59 = cur_rs2 == _GEN_134 & _T_17 ? _GEN_11 : _GEN_56; // @[forwading.scala 133:82]
  wire [63:0] _GEN_60 = cur_rs2 == _GEN_133 & _T_13 ? _GEN_6 : _GEN_57; // @[forwading.scala 126:82]
  wire  _GEN_61 = cur_rs2 == _GEN_133 & _T_13 ? _T_15 : _GEN_58; // @[forwading.scala 126:82]
  wire  _GEN_62 = cur_rs2 == _GEN_133 & _T_13 ? _GEN_8 : _GEN_59; // @[forwading.scala 126:82]
  wire [63:0] _GEN_63 = cur_rs2 == _GEN_132 & _T_9 ? _GEN_3 : _GEN_60; // @[forwading.scala 119:78]
  wire  _GEN_64 = cur_rs2 == _GEN_132 & _T_9 ? _T_11 : _GEN_61; // @[forwading.scala 119:78]
  wire  _GEN_65 = cur_rs2 == _GEN_132 & _T_9 ? _GEN_5 : _GEN_62; // @[forwading.scala 119:78]
  wire [63:0] _GEN_66 = cur_rs2 == _GEN_131 & _T_5 ? _GEN_0 : _GEN_63; // @[forwading.scala 112:78]
  wire  _GEN_67 = cur_rs2 == _GEN_131 & _T_5 ? _T_7 : _GEN_64; // @[forwading.scala 112:78]
  wire  _GEN_68 = cur_rs2 == _GEN_131 & _T_5 ? _GEN_2 : _GEN_65; // @[forwading.scala 112:78]
  wire  _GEN_69 = _T_1 & cur_rs2 == _GEN_130 | _GEN_68; // @[forwading.scala 110:60 forwading.scala 111:22]
  wire [63:0] _GEN_70 = _T_1 & cur_rs2 == _GEN_130 ? 64'h0 : _GEN_66; // @[forwading.scala 110:60 forwading.scala 58:62]
  wire  _GEN_71 = _T_1 & cur_rs2 == _GEN_130 ? 1'h0 : _GEN_67; // @[forwading.scala 110:60 forwading.scala 58:15]
  wire  _GEN_72 = cur_rs2 == 12'h0 ? 1'h0 : _GEN_69; // @[forwading.scala 108:30 forwading.scala 109:22]
  wire [63:0] _GEN_73 = cur_rs2 == 12'h0 ? 64'h0 : _GEN_70; // @[forwading.scala 108:30 forwading.scala 58:62]
  wire  _GEN_74 = cur_rs2 == 12'h0 ? 1'h0 : _GEN_71; // @[forwading.scala 108:30 forwading.scala 58:15]
  wire  rs2_wait = cur_rrs2 & _GEN_72; // @[forwading.scala 106:19 forwading.scala 58:41]
  wire  rs2_valid = cur_rrs2 & _GEN_74; // @[forwading.scala 106:19 forwading.scala 58:15]
  wire [63:0] _GEN_93 = hs_in ? io_id2df_rs1_d : rs1_d_r; // @[forwading.scala 150:16 forwading.scala 157:21 forwading.scala 30:30]
  wire [63:0] _GEN_96 = hs_in ? io_id2df_rs2_d : rs2_d_r; // @[forwading.scala 150:16 forwading.scala 160:21 forwading.scala 33:30]
  wire  _GEN_116 = (valid_r | state) & ~hs_out ? 1'h0 : io_id2df_valid; // @[forwading.scala 191:54 forwading.scala 189:20]
  wire  _GEN_117 = hs_out ? 1'h0 : valid_r; // @[forwading.scala 202:31 forwading.scala 203:25 forwading.scala 41:30]
  wire  _GEN_118 = hs_in | _GEN_117; // @[forwading.scala 200:30 forwading.scala 201:25]
  wire  _GEN_119 = hs_in & (rs1_wait | rs2_wait) | state; // @[forwading.scala 197:50 forwading.scala 198:23 forwading.scala 47:24]
  wire  _GEN_120 = hs_in & (rs1_wait | rs2_wait) ? 1'h0 : _GEN_118; // @[forwading.scala 197:50 forwading.scala 199:25]
  wire  _GEN_121 = ~state ? _GEN_119 : state; // @[forwading.scala 196:30 forwading.scala 47:24]
  wire  _GEN_122 = ~state ? _GEN_120 : valid_r; // @[forwading.scala 196:30 forwading.scala 41:30]
  wire  _GEN_123 = ~rs1_wait & ~rs2_wait ? 1'h0 : _GEN_121; // @[forwading.scala 207:43 forwading.scala 208:23]
  wire  _GEN_124 = ~rs1_wait & ~rs2_wait | _GEN_122; // @[forwading.scala 207:43 forwading.scala 209:25]
  wire  _GEN_125 = state ? _GEN_123 : _GEN_121; // @[forwading.scala 206:30]
  wire  _GEN_126 = state ? _GEN_124 : _GEN_122; // @[forwading.scala 206:30]
  wire  _GEN_128 = _io_id2df_stall_T & _GEN_125; // @[forwading.scala 190:25 forwading.scala 214:21]
  wire  _GEN_129 = _io_id2df_stall_T & _GEN_126; // @[forwading.scala 190:25 forwading.scala 215:21]
  assign io_id2df_drop = io_df2rr_drop; // @[forwading.scala 22:31]
  assign io_id2df_stall = io_df2rr_stall; // @[forwading.scala 23:52]
  assign io_id2df_ready = _io_id2df_stall_T & _GEN_116; // @[forwading.scala 190:25 forwading.scala 189:20]
  assign io_df2rr_inst = inst_r; // @[forwading.scala 217:25]
  assign io_df2rr_pc = pc_r; // @[forwading.scala 218:25]
  assign io_df2rr_excep_cause = excep_r_cause; // @[forwading.scala 219:25]
  assign io_df2rr_excep_tval = excep_r_tval; // @[forwading.scala 219:25]
  assign io_df2rr_excep_en = excep_r_en; // @[forwading.scala 219:25]
  assign io_df2rr_excep_pc = excep_r_pc; // @[forwading.scala 219:25]
  assign io_df2rr_excep_etype = excep_r_etype; // @[forwading.scala 219:25]
  assign io_df2rr_ctrl_aluOp = ctrl_r_aluOp; // @[forwading.scala 220:25]
  assign io_df2rr_ctrl_aluWidth = ctrl_r_aluWidth; // @[forwading.scala 220:25]
  assign io_df2rr_ctrl_dcMode = ctrl_r_dcMode; // @[forwading.scala 220:25]
  assign io_df2rr_ctrl_writeRegEn = ctrl_r_writeRegEn; // @[forwading.scala 220:25]
  assign io_df2rr_ctrl_writeCSREn = ctrl_r_writeCSREn; // @[forwading.scala 220:25]
  assign io_df2rr_ctrl_brType = ctrl_r_brType; // @[forwading.scala 220:25]
  assign io_df2rr_rs1 = rs1_r; // @[forwading.scala 221:25]
  assign io_df2rr_rrs1 = rrs1_r; // @[forwading.scala 222:25]
  assign io_df2rr_rs1_d = rs1_d_r; // @[forwading.scala 223:25]
  assign io_df2rr_rs2 = rs2_r; // @[forwading.scala 224:25]
  assign io_df2rr_rrs2 = rrs2_r; // @[forwading.scala 225:25]
  assign io_df2rr_rs2_d = rs2_d_r; // @[forwading.scala 226:25]
  assign io_df2rr_dst = dst_r; // @[forwading.scala 227:25]
  assign io_df2rr_dst_d = dst_d_r; // @[forwading.scala 228:25]
  assign io_df2rr_jmp_type = jmp_type_r; // @[forwading.scala 229:25]
  assign io_df2rr_special = special_r; // @[forwading.scala 230:25]
  assign io_df2rr_swap = swap_r; // @[forwading.scala 232:25]
  assign io_df2rr_indi = indi_r; // @[forwading.scala 231:25]
  assign io_df2rr_recov = recov_r; // @[forwading.scala 233:25]
  assign io_df2rr_valid = valid_r; // @[forwading.scala 234:25]
  always @(posedge clock) begin
    if (reset) begin // @[forwading.scala 24:30]
      inst_r <= 32'h0; // @[forwading.scala 24:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      inst_r <= io_id2df_inst; // @[forwading.scala 151:21]
    end
    if (reset) begin // @[forwading.scala 25:30]
      pc_r <= 64'h0; // @[forwading.scala 25:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      pc_r <= io_id2df_pc; // @[forwading.scala 152:21]
    end
    if (reset) begin // @[forwading.scala 26:30]
      excep_r_cause <= 64'h0; // @[forwading.scala 26:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      excep_r_cause <= io_id2df_excep_cause; // @[forwading.scala 153:21]
    end
    if (reset) begin // @[forwading.scala 26:30]
      excep_r_tval <= 64'h0; // @[forwading.scala 26:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      excep_r_tval <= io_id2df_excep_tval; // @[forwading.scala 153:21]
    end
    if (reset) begin // @[forwading.scala 26:30]
      excep_r_en <= 1'h0; // @[forwading.scala 26:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      excep_r_en <= io_id2df_excep_en; // @[forwading.scala 153:21]
    end
    if (reset) begin // @[forwading.scala 26:30]
      excep_r_pc <= 64'h0; // @[forwading.scala 26:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      excep_r_pc <= io_id2df_excep_pc; // @[forwading.scala 153:21]
    end
    if (reset) begin // @[forwading.scala 26:30]
      excep_r_etype <= 2'h0; // @[forwading.scala 26:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      excep_r_etype <= io_id2df_excep_etype; // @[forwading.scala 153:21]
    end
    if (reset) begin // @[forwading.scala 27:30]
      ctrl_r_aluOp <= 5'h0; // @[forwading.scala 27:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      ctrl_r_aluOp <= io_id2df_ctrl_aluOp; // @[forwading.scala 154:21]
    end
    if (reset) begin // @[forwading.scala 27:30]
      ctrl_r_aluWidth <= 1'h0; // @[forwading.scala 27:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      ctrl_r_aluWidth <= io_id2df_ctrl_aluWidth; // @[forwading.scala 154:21]
    end
    if (reset) begin // @[forwading.scala 27:30]
      ctrl_r_dcMode <= 5'h0; // @[forwading.scala 27:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      ctrl_r_dcMode <= io_id2df_ctrl_dcMode; // @[forwading.scala 154:21]
    end
    if (reset) begin // @[forwading.scala 27:30]
      ctrl_r_writeRegEn <= 1'h0; // @[forwading.scala 27:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      ctrl_r_writeRegEn <= io_id2df_ctrl_writeRegEn; // @[forwading.scala 154:21]
    end
    if (reset) begin // @[forwading.scala 27:30]
      ctrl_r_writeCSREn <= 1'h0; // @[forwading.scala 27:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      ctrl_r_writeCSREn <= io_id2df_ctrl_writeCSREn; // @[forwading.scala 154:21]
    end
    if (reset) begin // @[forwading.scala 27:30]
      ctrl_r_brType <= 3'h0; // @[forwading.scala 27:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      ctrl_r_brType <= io_id2df_ctrl_brType; // @[forwading.scala 154:21]
    end
    if (reset) begin // @[forwading.scala 28:30]
      rs1_r <= 5'h0; // @[forwading.scala 28:30]
    end else if (hs_in) begin // @[forwading.scala 59:26]
      rs1_r <= io_id2df_rs1;
    end
    if (reset) begin // @[forwading.scala 29:30]
      rrs1_r <= 1'h0; // @[forwading.scala 29:30]
    end else if (hs_in | state) begin // @[forwading.scala 170:37]
      if (rs1_valid & cur_rrs1) begin // @[forwading.scala 171:36]
        rrs1_r <= 1'h0; // @[forwading.scala 172:21]
      end else begin
        rrs1_r <= cur_rrs1;
      end
    end else begin
      rrs1_r <= cur_rrs1;
    end
    if (reset) begin // @[forwading.scala 30:30]
      rs1_d_r <= 64'h0; // @[forwading.scala 30:30]
    end else if (hs_in | state) begin // @[forwading.scala 170:37]
      if (rs1_valid & cur_rrs1) begin // @[forwading.scala 171:36]
        if (cur_rrs1) begin // @[forwading.scala 63:19]
          rs1_d_r <= _GEN_34;
        end else begin
          rs1_d_r <= 64'h0; // @[forwading.scala 57:62]
        end
      end else begin
        rs1_d_r <= _GEN_93;
      end
    end else begin
      rs1_d_r <= _GEN_93;
    end
    if (reset) begin // @[forwading.scala 31:30]
      rs2_r <= 12'h0; // @[forwading.scala 31:30]
    end else if (hs_in) begin // @[forwading.scala 61:26]
      rs2_r <= io_id2df_rs2;
    end
    if (reset) begin // @[forwading.scala 32:30]
      rrs2_r <= 1'h0; // @[forwading.scala 32:30]
    end else if (hs_in | state) begin // @[forwading.scala 170:37]
      if (rs2_valid & cur_rrs2) begin // @[forwading.scala 175:36]
        rrs2_r <= 1'h0; // @[forwading.scala 176:21]
      end else begin
        rrs2_r <= cur_rrs2;
      end
    end else begin
      rrs2_r <= cur_rrs2;
    end
    if (reset) begin // @[forwading.scala 33:30]
      rs2_d_r <= 64'h0; // @[forwading.scala 33:30]
    end else if (hs_in | state) begin // @[forwading.scala 170:37]
      if (rs2_valid & cur_rrs2) begin // @[forwading.scala 175:36]
        if (cur_rrs2) begin // @[forwading.scala 106:19]
          rs2_d_r <= _GEN_73;
        end else begin
          rs2_d_r <= 64'h0; // @[forwading.scala 58:62]
        end
      end else begin
        rs2_d_r <= _GEN_96;
      end
    end else begin
      rs2_d_r <= _GEN_96;
    end
    if (reset) begin // @[forwading.scala 34:30]
      dst_r <= 5'h0; // @[forwading.scala 34:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      dst_r <= io_id2df_dst; // @[forwading.scala 161:21]
    end
    if (reset) begin // @[forwading.scala 35:30]
      dst_d_r <= 64'h0; // @[forwading.scala 35:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      dst_d_r <= io_id2df_dst_d; // @[forwading.scala 162:21]
    end
    if (reset) begin // @[forwading.scala 36:30]
      jmp_type_r <= 2'h0; // @[forwading.scala 36:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      jmp_type_r <= io_id2df_jmp_type; // @[forwading.scala 163:21]
    end
    if (reset) begin // @[forwading.scala 37:30]
      special_r <= 2'h0; // @[forwading.scala 37:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      special_r <= io_id2df_special; // @[forwading.scala 164:21]
    end
    if (reset) begin // @[forwading.scala 38:30]
      indi_r <= 2'h0; // @[forwading.scala 38:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      indi_r <= io_id2df_indi; // @[forwading.scala 165:21]
    end
    if (reset) begin // @[forwading.scala 39:30]
      swap_r <= 6'h0; // @[forwading.scala 39:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      swap_r <= io_id2df_swap; // @[forwading.scala 166:21]
    end
    if (reset) begin // @[forwading.scala 40:30]
      recov_r <= 1'h0; // @[forwading.scala 40:30]
    end else if (hs_in) begin // @[forwading.scala 150:16]
      recov_r <= io_id2df_recov; // @[forwading.scala 167:21]
    end
    if (reset) begin // @[forwading.scala 41:30]
      valid_r <= 1'h0; // @[forwading.scala 41:30]
    end else begin
      valid_r <= _GEN_129;
    end
    if (reset) begin // @[forwading.scala 43:30]
      pre_dst <= 5'h0; // @[forwading.scala 43:30]
    end else if (hs_in) begin // @[forwading.scala 181:16]
      pre_dst <= io_id2df_dst; // @[forwading.scala 182:17]
    end
    if (reset) begin // @[forwading.scala 44:30]
      pre_wr <= 1'h0; // @[forwading.scala 44:30]
    end else if (hs_in) begin // @[forwading.scala 181:16]
      pre_wr <= io_id2df_ctrl_writeRegEn; // @[forwading.scala 183:17]
    end else if (hs_out) begin // @[forwading.scala 184:23]
      pre_wr <= 1'h0; // @[forwading.scala 185:17]
    end
    if (reset) begin // @[forwading.scala 47:24]
      state <= 1'h0; // @[forwading.scala 47:24]
    end else begin
      state <= _GEN_128;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inst_r = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  pc_r = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  excep_r_cause = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  excep_r_tval = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  excep_r_en = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  excep_r_pc = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  excep_r_etype = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  ctrl_r_aluOp = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  ctrl_r_aluWidth = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  ctrl_r_dcMode = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  ctrl_r_writeRegEn = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ctrl_r_writeCSREn = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ctrl_r_brType = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  rs1_r = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  rrs1_r = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  rs1_d_r = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  rs2_r = _RAND_16[11:0];
  _RAND_17 = {1{`RANDOM}};
  rrs2_r = _RAND_17[0:0];
  _RAND_18 = {2{`RANDOM}};
  rs2_d_r = _RAND_18[63:0];
  _RAND_19 = {1{`RANDOM}};
  dst_r = _RAND_19[4:0];
  _RAND_20 = {2{`RANDOM}};
  dst_d_r = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  jmp_type_r = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  special_r = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  indi_r = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  swap_r = _RAND_24[5:0];
  _RAND_25 = {1{`RANDOM}};
  recov_r = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_r = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  pre_dst = _RAND_27[4:0];
  _RAND_28 = {1{`RANDOM}};
  pre_wr = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  state = _RAND_29[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_ReadRegs(
  input         clock,
  input         reset,
  input  [31:0] io_df2rr_inst,
  input  [63:0] io_df2rr_pc,
  input  [63:0] io_df2rr_excep_cause,
  input  [63:0] io_df2rr_excep_tval,
  input         io_df2rr_excep_en,
  input  [63:0] io_df2rr_excep_pc,
  input  [1:0]  io_df2rr_excep_etype,
  input  [4:0]  io_df2rr_ctrl_aluOp,
  input         io_df2rr_ctrl_aluWidth,
  input  [4:0]  io_df2rr_ctrl_dcMode,
  input         io_df2rr_ctrl_writeRegEn,
  input         io_df2rr_ctrl_writeCSREn,
  input  [2:0]  io_df2rr_ctrl_brType,
  input  [4:0]  io_df2rr_rs1,
  input         io_df2rr_rrs1,
  input  [63:0] io_df2rr_rs1_d,
  input  [11:0] io_df2rr_rs2,
  input         io_df2rr_rrs2,
  input  [63:0] io_df2rr_rs2_d,
  input  [4:0]  io_df2rr_dst,
  input  [63:0] io_df2rr_dst_d,
  input  [1:0]  io_df2rr_jmp_type,
  input  [1:0]  io_df2rr_special,
  input  [5:0]  io_df2rr_swap,
  input  [1:0]  io_df2rr_indi,
  output        io_df2rr_drop,
  output        io_df2rr_stall,
  input         io_df2rr_recov,
  input         io_df2rr_valid,
  output        io_df2rr_ready,
  output [31:0] io_rr2ex_inst,
  output [63:0] io_rr2ex_pc,
  output [63:0] io_rr2ex_excep_cause,
  output [63:0] io_rr2ex_excep_tval,
  output        io_rr2ex_excep_en,
  output [63:0] io_rr2ex_excep_pc,
  output [1:0]  io_rr2ex_excep_etype,
  output [4:0]  io_rr2ex_ctrl_aluOp,
  output        io_rr2ex_ctrl_aluWidth,
  output [4:0]  io_rr2ex_ctrl_dcMode,
  output        io_rr2ex_ctrl_writeRegEn,
  output        io_rr2ex_ctrl_writeCSREn,
  output [2:0]  io_rr2ex_ctrl_brType,
  output [63:0] io_rr2ex_rs1_d,
  output [11:0] io_rr2ex_rs2,
  output [63:0] io_rr2ex_rs2_d,
  output [4:0]  io_rr2ex_dst,
  output [63:0] io_rr2ex_dst_d,
  output [11:0] io_rr2ex_rcsr_id,
  output [1:0]  io_rr2ex_jmp_type,
  output [1:0]  io_rr2ex_special,
  output [1:0]  io_rr2ex_indi,
  input         io_rr2ex_drop,
  input         io_rr2ex_stall,
  output        io_rr2ex_recov,
  output        io_rr2ex_valid,
  input         io_rr2ex_ready,
  output [4:0]  io_rs1Read_id,
  input  [63:0] io_rs1Read_data,
  output [4:0]  io_rs2Read_id,
  input  [63:0] io_rs2Read_data,
  output [11:0] io_csrRead_id,
  input  [63:0] io_csrRead_data,
  input         io_csrRead_is_err,
  output [4:0]  io_d_rr_id,
  output [63:0] io_d_rr_data,
  output [1:0]  io_d_rr_state
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
`endif // RANDOMIZE_REG_INIT
  reg  drop_r; // @[readregs.scala 18:30]
  reg  stall_r; // @[readregs.scala 20:30]
  reg  recov_r; // @[readregs.scala 22:30]
  wire  drop_in = io_rr2ex_drop | drop_r; // @[readregs.scala 26:37]
  wire  _io_df2rr_stall_T = ~io_rr2ex_drop; // @[readregs.scala 28:36]
  reg [31:0] inst_r; // @[readregs.scala 29:30]
  reg [63:0] pc_r; // @[readregs.scala 30:30]
  reg [63:0] excep_r_cause; // @[readregs.scala 31:30]
  reg [63:0] excep_r_tval; // @[readregs.scala 31:30]
  reg  excep_r_en; // @[readregs.scala 31:30]
  reg [63:0] excep_r_pc; // @[readregs.scala 31:30]
  reg [1:0] excep_r_etype; // @[readregs.scala 31:30]
  reg [4:0] ctrl_r_aluOp; // @[readregs.scala 32:30]
  reg  ctrl_r_aluWidth; // @[readregs.scala 32:30]
  reg [4:0] ctrl_r_dcMode; // @[readregs.scala 32:30]
  reg  ctrl_r_writeRegEn; // @[readregs.scala 32:30]
  reg  ctrl_r_writeCSREn; // @[readregs.scala 32:30]
  reg [2:0] ctrl_r_brType; // @[readregs.scala 32:30]
  reg [63:0] rs1_d_r; // @[readregs.scala 34:30]
  reg [11:0] rs2_r; // @[readregs.scala 35:30]
  reg [63:0] rs2_d_r; // @[readregs.scala 36:30]
  reg [4:0] dst_r; // @[readregs.scala 37:30]
  reg [63:0] dst_d_r; // @[readregs.scala 38:30]
  reg [11:0] rcsr_id_r; // @[readregs.scala 39:30]
  reg [1:0] jmp_type_r; // @[readregs.scala 40:30]
  reg [1:0] special_r; // @[readregs.scala 41:30]
  reg [1:0] indi_r; // @[readregs.scala 42:30]
  reg  valid_r; // @[readregs.scala 44:30]
  wire  hs_in = io_df2rr_ready & io_df2rr_valid; // @[readregs.scala 46:34]
  wire  hs_out = io_rr2ex_ready & io_rr2ex_valid; // @[readregs.scala 47:34]
  wire [63:0] rs1_bef = io_df2rr_rrs1 ? io_rs1Read_data : io_df2rr_rs1_d; // @[readregs.scala 52:22]
  wire [63:0] _rs2_bef_T_2 = io_df2rr_rrs2 ? io_rs2Read_data : io_df2rr_rs2_d; // @[readregs.scala 53:98]
  wire [63:0] rs2_bef = io_df2rr_ctrl_writeCSREn | io_df2rr_excep_en ? io_csrRead_data : _rs2_bef_T_2; // @[readregs.scala 53:22]
  wire [63:0] _rs1_d_r_T_2 = 2'h1 == io_df2rr_swap[5:4] ? rs1_bef : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _rs2_d_r_T_2 = 2'h1 == io_df2rr_swap[3:2] ? rs1_bef : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _dst_d_r_T_2 = 2'h1 == io_df2rr_swap[1:0] ? rs1_bef : 64'h0; // @[Mux.scala 80:57]
  wire  _T = io_df2rr_ctrl_writeCSREn & io_csrRead_is_err; // @[readregs.scala 78:39]
  wire  _GEN_2 = io_df2rr_ctrl_writeCSREn & io_csrRead_is_err | io_df2rr_excep_en; // @[readregs.scala 78:60 readregs.scala 81:29 readregs.scala 65:21]
  wire  _GEN_6 = io_df2rr_ctrl_writeCSREn & io_csrRead_is_err | io_df2rr_recov; // @[readregs.scala 78:60 readregs.scala 24:57 readregs.scala 77:21]
  wire  _GEN_39 = hs_in & _T; // @[readregs.scala 62:16 readregs.scala 19:21]
  wire  _GEN_41 = valid_r & ~hs_out ? 1'h0 : io_df2rr_valid; // @[readregs.scala 92:33 readregs.scala 90:20]
  wire  _GEN_43 = hs_out ? 1'h0 : valid_r; // @[readregs.scala 100:27 readregs.scala 101:21 readregs.scala 44:30]
  wire  _GEN_44 = hs_in | _GEN_43; // @[readregs.scala 98:20 readregs.scala 99:21]
  wire  _GEN_45 = _io_df2rr_stall_T & _GEN_44; // @[readregs.scala 97:25 readregs.scala 104:17]
  assign io_df2rr_drop = io_rr2ex_drop | drop_r; // @[readregs.scala 26:37]
  assign io_df2rr_stall = stall_r & ~io_rr2ex_drop | io_rr2ex_stall; // @[readregs.scala 28:52]
  assign io_df2rr_ready = ~drop_in & _GEN_41; // @[readregs.scala 91:19 readregs.scala 90:20]
  assign io_rr2ex_inst = inst_r; // @[readregs.scala 106:25]
  assign io_rr2ex_pc = pc_r; // @[readregs.scala 107:25]
  assign io_rr2ex_excep_cause = excep_r_cause; // @[readregs.scala 108:25]
  assign io_rr2ex_excep_tval = excep_r_tval; // @[readregs.scala 108:25]
  assign io_rr2ex_excep_en = excep_r_en; // @[readregs.scala 108:25]
  assign io_rr2ex_excep_pc = excep_r_pc; // @[readregs.scala 108:25]
  assign io_rr2ex_excep_etype = excep_r_etype; // @[readregs.scala 108:25]
  assign io_rr2ex_ctrl_aluOp = ctrl_r_aluOp; // @[readregs.scala 109:25]
  assign io_rr2ex_ctrl_aluWidth = ctrl_r_aluWidth; // @[readregs.scala 109:25]
  assign io_rr2ex_ctrl_dcMode = ctrl_r_dcMode; // @[readregs.scala 109:25]
  assign io_rr2ex_ctrl_writeRegEn = ctrl_r_writeRegEn; // @[readregs.scala 109:25]
  assign io_rr2ex_ctrl_writeCSREn = ctrl_r_writeCSREn; // @[readregs.scala 109:25]
  assign io_rr2ex_ctrl_brType = ctrl_r_brType; // @[readregs.scala 109:25]
  assign io_rr2ex_rs1_d = rs1_d_r; // @[readregs.scala 111:25]
  assign io_rr2ex_rs2 = rs2_r; // @[readregs.scala 112:25]
  assign io_rr2ex_rs2_d = rs2_d_r; // @[readregs.scala 113:25]
  assign io_rr2ex_dst = dst_r; // @[readregs.scala 114:25]
  assign io_rr2ex_dst_d = dst_d_r; // @[readregs.scala 115:25]
  assign io_rr2ex_rcsr_id = rcsr_id_r; // @[readregs.scala 116:25]
  assign io_rr2ex_jmp_type = jmp_type_r; // @[readregs.scala 117:25]
  assign io_rr2ex_special = special_r; // @[readregs.scala 118:25]
  assign io_rr2ex_indi = indi_r; // @[readregs.scala 119:25]
  assign io_rr2ex_recov = recov_r; // @[readregs.scala 120:25]
  assign io_rr2ex_valid = valid_r; // @[readregs.scala 121:25]
  assign io_rs1Read_id = io_df2rr_rs1; // @[readregs.scala 49:19]
  assign io_rs2Read_id = io_df2rr_rs2[4:0]; // @[readregs.scala 50:34]
  assign io_csrRead_id = io_df2rr_rs2; // @[readregs.scala 51:19]
  assign io_d_rr_id = dst_r; // @[readregs.scala 123:21]
  assign io_d_rr_data = dst_d_r; // @[readregs.scala 124:21]
  assign io_d_rr_state = valid_r ? 2'h2 : 2'h0; // @[readregs.scala 125:27]
  always @(posedge clock) begin
    if (reset) begin // @[readregs.scala 18:30]
      drop_r <= 1'h0; // @[readregs.scala 18:30]
    end else begin
      drop_r <= _GEN_39;
    end
    if (reset) begin // @[readregs.scala 20:30]
      stall_r <= 1'h0; // @[readregs.scala 20:30]
    end else begin
      stall_r <= _GEN_39;
    end
    if (reset) begin // @[readregs.scala 22:30]
      recov_r <= 1'h0; // @[readregs.scala 22:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      recov_r <= _GEN_6;
    end
    if (reset) begin // @[readregs.scala 29:30]
      inst_r <= 32'h0; // @[readregs.scala 29:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      inst_r <= io_df2rr_inst; // @[readregs.scala 63:21]
    end
    if (reset) begin // @[readregs.scala 30:30]
      pc_r <= 64'h0; // @[readregs.scala 30:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      pc_r <= io_df2rr_pc; // @[readregs.scala 64:21]
    end
    if (reset) begin // @[readregs.scala 31:30]
      excep_r_cause <= 64'h0; // @[readregs.scala 31:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[readregs.scala 78:60]
        excep_r_cause <= 64'h2; // @[readregs.scala 79:29]
      end else begin
        excep_r_cause <= io_df2rr_excep_cause; // @[readregs.scala 65:21]
      end
    end
    if (reset) begin // @[readregs.scala 31:30]
      excep_r_tval <= 64'h0; // @[readregs.scala 31:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[readregs.scala 78:60]
        excep_r_tval <= {{32'd0}, io_df2rr_inst}; // @[readregs.scala 80:29]
      end else begin
        excep_r_tval <= io_df2rr_excep_tval; // @[readregs.scala 65:21]
      end
    end
    if (reset) begin // @[readregs.scala 31:30]
      excep_r_en <= 1'h0; // @[readregs.scala 31:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      excep_r_en <= _GEN_2;
    end
    if (reset) begin // @[readregs.scala 31:30]
      excep_r_pc <= 64'h0; // @[readregs.scala 31:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[readregs.scala 78:60]
        excep_r_pc <= io_df2rr_pc; // @[readregs.scala 82:29]
      end else begin
        excep_r_pc <= io_df2rr_excep_pc; // @[readregs.scala 65:21]
      end
    end
    if (reset) begin // @[readregs.scala 31:30]
      excep_r_etype <= 2'h0; // @[readregs.scala 31:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[readregs.scala 78:60]
        excep_r_etype <= 2'h0; // @[readregs.scala 83:29]
      end else begin
        excep_r_etype <= io_df2rr_excep_etype; // @[readregs.scala 65:21]
      end
    end
    if (reset) begin // @[readregs.scala 32:30]
      ctrl_r_aluOp <= 5'h0; // @[readregs.scala 32:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[readregs.scala 78:60]
        ctrl_r_aluOp <= 5'h0; // @[readregs.scala 85:25]
      end else begin
        ctrl_r_aluOp <= io_df2rr_ctrl_aluOp; // @[readregs.scala 66:21]
      end
    end
    if (reset) begin // @[readregs.scala 32:30]
      ctrl_r_aluWidth <= 1'h0; // @[readregs.scala 32:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[readregs.scala 78:60]
        ctrl_r_aluWidth <= 1'h0; // @[readregs.scala 85:25]
      end else begin
        ctrl_r_aluWidth <= io_df2rr_ctrl_aluWidth; // @[readregs.scala 66:21]
      end
    end
    if (reset) begin // @[readregs.scala 32:30]
      ctrl_r_dcMode <= 5'h0; // @[readregs.scala 32:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[readregs.scala 78:60]
        ctrl_r_dcMode <= 5'h0; // @[readregs.scala 85:25]
      end else begin
        ctrl_r_dcMode <= io_df2rr_ctrl_dcMode; // @[readregs.scala 66:21]
      end
    end
    if (reset) begin // @[readregs.scala 32:30]
      ctrl_r_writeRegEn <= 1'h0; // @[readregs.scala 32:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[readregs.scala 78:60]
        ctrl_r_writeRegEn <= 1'h0; // @[readregs.scala 85:25]
      end else begin
        ctrl_r_writeRegEn <= io_df2rr_ctrl_writeRegEn; // @[readregs.scala 66:21]
      end
    end
    if (reset) begin // @[readregs.scala 32:30]
      ctrl_r_writeCSREn <= 1'h0; // @[readregs.scala 32:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[readregs.scala 78:60]
        ctrl_r_writeCSREn <= 1'h0; // @[readregs.scala 85:25]
      end else begin
        ctrl_r_writeCSREn <= io_df2rr_ctrl_writeCSREn; // @[readregs.scala 66:21]
      end
    end
    if (reset) begin // @[readregs.scala 32:30]
      ctrl_r_brType <= 3'h0; // @[readregs.scala 32:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[readregs.scala 78:60]
        ctrl_r_brType <= 3'h0; // @[readregs.scala 85:25]
      end else begin
        ctrl_r_brType <= io_df2rr_ctrl_brType; // @[readregs.scala 66:21]
      end
    end
    if (reset) begin // @[readregs.scala 34:30]
      rs1_d_r <= 64'h0; // @[readregs.scala 34:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      if (2'h3 == io_df2rr_swap[5:4]) begin // @[Mux.scala 80:57]
        rs1_d_r <= io_df2rr_dst_d;
      end else if (2'h2 == io_df2rr_swap[5:4]) begin // @[Mux.scala 80:57]
        rs1_d_r <= rs2_bef;
      end else begin
        rs1_d_r <= _rs1_d_r_T_2;
      end
    end
    if (reset) begin // @[readregs.scala 35:30]
      rs2_r <= 12'h0; // @[readregs.scala 35:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      rs2_r <= io_df2rr_rs2; // @[readregs.scala 69:21]
    end
    if (reset) begin // @[readregs.scala 36:30]
      rs2_d_r <= 64'h0; // @[readregs.scala 36:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      if (2'h3 == io_df2rr_swap[3:2]) begin // @[Mux.scala 80:57]
        rs2_d_r <= io_df2rr_dst_d;
      end else if (2'h2 == io_df2rr_swap[3:2]) begin // @[Mux.scala 80:57]
        rs2_d_r <= rs2_bef;
      end else begin
        rs2_d_r <= _rs2_d_r_T_2;
      end
    end
    if (reset) begin // @[readregs.scala 37:30]
      dst_r <= 5'h0; // @[readregs.scala 37:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      dst_r <= io_df2rr_dst; // @[readregs.scala 71:21]
    end
    if (reset) begin // @[readregs.scala 38:30]
      dst_d_r <= 64'h0; // @[readregs.scala 38:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      if (2'h3 == io_df2rr_swap[1:0]) begin // @[Mux.scala 80:57]
        dst_d_r <= io_df2rr_dst_d;
      end else if (2'h2 == io_df2rr_swap[1:0]) begin // @[Mux.scala 80:57]
        dst_d_r <= rs2_bef;
      end else begin
        dst_d_r <= _dst_d_r_T_2;
      end
    end
    if (reset) begin // @[readregs.scala 39:30]
      rcsr_id_r <= 12'h0; // @[readregs.scala 39:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn) begin // @[readregs.scala 73:27]
        rcsr_id_r <= io_df2rr_rs2;
      end else begin
        rcsr_id_r <= 12'h0;
      end
    end
    if (reset) begin // @[readregs.scala 40:30]
      jmp_type_r <= 2'h0; // @[readregs.scala 40:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[readregs.scala 78:60]
        jmp_type_r <= 2'h0; // @[readregs.scala 86:25]
      end else begin
        jmp_type_r <= io_df2rr_jmp_type; // @[readregs.scala 74:21]
      end
    end
    if (reset) begin // @[readregs.scala 41:30]
      special_r <= 2'h0; // @[readregs.scala 41:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[readregs.scala 78:60]
        special_r <= 2'h0; // @[readregs.scala 87:25]
      end else begin
        special_r <= io_df2rr_special; // @[readregs.scala 75:21]
      end
    end
    if (reset) begin // @[readregs.scala 42:30]
      indi_r <= 2'h0; // @[readregs.scala 42:30]
    end else if (hs_in) begin // @[readregs.scala 62:16]
      indi_r <= io_df2rr_indi; // @[readregs.scala 76:21]
    end
    if (reset) begin // @[readregs.scala 44:30]
      valid_r <= 1'h0; // @[readregs.scala 44:30]
    end else begin
      valid_r <= _GEN_45;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  drop_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  stall_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  recov_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  inst_r = _RAND_3[31:0];
  _RAND_4 = {2{`RANDOM}};
  pc_r = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  excep_r_cause = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  excep_r_tval = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  excep_r_en = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  excep_r_pc = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  excep_r_etype = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  ctrl_r_aluOp = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  ctrl_r_aluWidth = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ctrl_r_dcMode = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  ctrl_r_writeRegEn = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  ctrl_r_writeCSREn = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  ctrl_r_brType = _RAND_15[2:0];
  _RAND_16 = {2{`RANDOM}};
  rs1_d_r = _RAND_16[63:0];
  _RAND_17 = {1{`RANDOM}};
  rs2_r = _RAND_17[11:0];
  _RAND_18 = {2{`RANDOM}};
  rs2_d_r = _RAND_18[63:0];
  _RAND_19 = {1{`RANDOM}};
  dst_r = _RAND_19[4:0];
  _RAND_20 = {2{`RANDOM}};
  dst_d_r = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  rcsr_id_r = _RAND_21[11:0];
  _RAND_22 = {1{`RANDOM}};
  jmp_type_r = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  special_r = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  indi_r = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  valid_r = _RAND_25[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_MUL(
  input         clock,
  input         reset,
  input  [63:0] io_a,
  input  [63:0] io_b,
  input  [4:0]  io_aluop,
  input         io_en,
  output [63:0] io_out,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] out_r; // @[muldiv.scala 20:30]
  reg [63:0] val1; // @[muldiv.scala 21:30]
  reg [63:0] val2; // @[muldiv.scala 22:30]
  reg [4:0] aluop_r; // @[muldiv.scala 23:33]
  reg  valid_r; // @[muldiv.scala 24:30]
  reg [1:0] state; // @[muldiv.scala 26:24]
  wire  _T = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire [127:0] _out_r_T = val1 * val2; // @[muldiv.scala 42:34]
  wire [127:0] _out_r_T_4 = $signed(val1) * $signed(val2); // @[muldiv.scala 43:42]
  wire [64:0] _out_r_T_9 = {1'b0,$signed(val2)}; // @[muldiv.scala 45:41]
  wire [128:0] _out_r_T_10 = $signed(val1) * $signed(_out_r_T_9); // @[muldiv.scala 45:41]
  wire [127:0] _out_r_T_12 = _out_r_T_10[127:0]; // @[muldiv.scala 45:41]
  wire [63:0] _out_r_T_15 = _out_r_T_12[127:64]; // @[muldiv.scala 45:65]
  wire [63:0] _out_r_T_17 = 5'hd == aluop_r ? _out_r_T[63:0] : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _out_r_T_19 = 5'he == aluop_r ? _out_r_T_4[127:64] : _out_r_T_17; // @[Mux.scala 80:57]
  wire [63:0] _out_r_T_21 = 5'hf == aluop_r ? _out_r_T[127:64] : _out_r_T_19; // @[Mux.scala 80:57]
  wire  _GEN_5 = _T_1 | valid_r; // @[Conditional.scala 39:67 muldiv.scala 47:21 muldiv.scala 24:30]
  assign io_out = out_r; // @[muldiv.scala 28:12]
  assign io_valid = valid_r; // @[muldiv.scala 29:14]
  always @(posedge clock) begin
    if (reset) begin // @[muldiv.scala 20:30]
      out_r <= 64'h0; // @[muldiv.scala 20:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (5'h10 == aluop_r) begin // @[Mux.scala 80:57]
          out_r <= _out_r_T_15;
        end else begin
          out_r <= _out_r_T_21;
        end
      end
    end
    if (reset) begin // @[muldiv.scala 21:30]
      val1 <= 64'h0; // @[muldiv.scala 21:30]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_en) begin // @[muldiv.scala 33:24]
        val1 <= io_a; // @[muldiv.scala 35:22]
      end
    end
    if (reset) begin // @[muldiv.scala 22:30]
      val2 <= 64'h0; // @[muldiv.scala 22:30]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_en) begin // @[muldiv.scala 33:24]
        val2 <= io_b; // @[muldiv.scala 36:22]
      end
    end
    if (reset) begin // @[muldiv.scala 23:33]
      aluop_r <= 5'h0; // @[muldiv.scala 23:33]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_en) begin // @[muldiv.scala 33:24]
        aluop_r <= io_aluop; // @[muldiv.scala 37:25]
      end
    end
    if (reset) begin // @[muldiv.scala 24:30]
      valid_r <= 1'h0; // @[muldiv.scala 24:30]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_r <= 1'h0; // @[muldiv.scala 32:21]
    end else begin
      valid_r <= _GEN_5;
    end
    if (reset) begin // @[muldiv.scala 26:24]
      state <= 2'h0; // @[muldiv.scala 26:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_en) begin // @[muldiv.scala 33:24]
        state <= 2'h1; // @[muldiv.scala 34:23]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      state <= 2'h0; // @[muldiv.scala 48:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  out_r = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  val1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  val2 = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  aluop_r = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_DIV(
  input         clock,
  input         reset,
  input         io_alu64,
  input  [63:0] io_a,
  input  [63:0] io_b,
  input         io_sign,
  input         io_en,
  output [63:0] io_qua,
  output [63:0] io_rem,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] quatient; // @[muldiv.scala 67:27]
  reg [127:0] val1; // @[muldiv.scala 68:26]
  reg [127:0] val2; // @[muldiv.scala 69:26]
  reg  qua_sign; // @[muldiv.scala 70:27]
  reg  rem_sign; // @[muldiv.scala 71:27]
  reg [6:0] iter; // @[muldiv.scala 72:26]
  reg  pre_alu64; // @[muldiv.scala 73:28]
  reg [1:0] state; // @[muldiv.scala 75:24]
  wire  _T = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _val1_T_2 = io_sign & io_a[63]; // @[muldiv.scala 84:61]
  wire [63:0] _val1_T_3 = ~io_a; // @[muldiv.scala 84:82]
  wire [63:0] _val1_T_5 = _val1_T_3 + 64'h1; // @[muldiv.scala 84:87]
  wire [63:0] val1_lo = io_sign & io_a[63] ? _val1_T_5 : io_a; // @[muldiv.scala 84:52]
  wire [127:0] _val1_T_6 = {64'h0,val1_lo}; // @[Cat.scala 30:58]
  wire [63:0] _val2_T_3 = ~io_b; // @[muldiv.scala 85:62]
  wire [63:0] _val2_T_5 = _val2_T_3 + 64'h1; // @[muldiv.scala 85:67]
  wire [63:0] val2_hi = io_sign & io_b[63] ? _val2_T_5 : io_b; // @[muldiv.scala 85:32]
  wire [127:0] _val2_T_6 = {val2_hi,64'h0}; // @[Cat.scala 30:58]
  wire  _T_1 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire [6:0] _iter_T_1 = iter + 7'h1; // @[muldiv.scala 95:30]
  wire [62:0] quatient_hi = quatient[62:0]; // @[muldiv.scala 97:45]
  wire [63:0] _quatient_T = {quatient_hi,1'h1}; // @[Cat.scala 30:58]
  wire [127:0] _val1_T_8 = val1 - val2; // @[muldiv.scala 98:34]
  wire [127:0] _val2_T_7 = {{1'd0}, val2[127:1]}; // @[muldiv.scala 99:34]
  wire [63:0] _quatient_T_1 = {quatient_hi,1'h0}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_8 = val1 >= val2 ? _quatient_T : _quatient_T_1; // @[muldiv.scala 96:35 muldiv.scala 97:30 muldiv.scala 101:30]
  wire [127:0] _GEN_9 = val1 >= val2 ? _val1_T_8 : val1; // @[muldiv.scala 96:35 muldiv.scala 98:26 muldiv.scala 68:26]
  wire [127:0] _GEN_10 = val1 >= val2 ? _val2_T_7 : _val2_T_7; // @[muldiv.scala 96:35 muldiv.scala 99:26 muldiv.scala 102:26]
  wire [63:0] _sign_qua_T = ~quatient; // @[muldiv.scala 107:46]
  wire [63:0] _sign_qua_T_2 = _sign_qua_T + 64'h1; // @[muldiv.scala 107:56]
  wire [63:0] sign_qua = qua_sign ? _sign_qua_T_2 : quatient; // @[muldiv.scala 107:35]
  wire [63:0] _sign_rem_T_1 = ~val1[63:0]; // @[muldiv.scala 108:46]
  wire [63:0] _sign_rem_T_3 = _sign_rem_T_1 + 64'h1; // @[muldiv.scala 108:58]
  wire [63:0] sign_rem = rem_sign ? _sign_rem_T_3 : val1[63:0]; // @[muldiv.scala 108:35]
  wire [31:0] io_qua_hi = sign_qua[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] io_qua_lo = sign_qua[31:0]; // @[muldiv.scala 109:90]
  wire [63:0] _io_qua_T_2 = {io_qua_hi,io_qua_lo}; // @[Cat.scala 30:58]
  wire [63:0] _io_qua_T_3 = pre_alu64 ? sign_qua : _io_qua_T_2; // @[muldiv.scala 109:32]
  wire [31:0] io_rem_hi = sign_rem[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] io_rem_lo = sign_rem[31:0]; // @[muldiv.scala 110:90]
  wire [63:0] _io_rem_T_2 = {io_rem_hi,io_rem_lo}; // @[Cat.scala 30:58]
  wire [63:0] _io_rem_T_3 = pre_alu64 ? sign_rem : _io_rem_T_2; // @[muldiv.scala 110:32]
  wire  _GEN_16 = iter <= 7'h40 ? 1'h0 : 1'h1; // @[muldiv.scala 94:39 muldiv.scala 79:14 muldiv.scala 106:26]
  wire [63:0] _GEN_17 = iter <= 7'h40 ? 64'h0 : _io_qua_T_3; // @[muldiv.scala 94:39 muldiv.scala 77:12 muldiv.scala 109:26]
  wire [63:0] _GEN_18 = iter <= 7'h40 ? 64'h0 : _io_rem_T_3; // @[muldiv.scala 94:39 muldiv.scala 78:12 muldiv.scala 110:26]
  wire  _GEN_24 = _T_1 & _GEN_16; // @[Conditional.scala 39:67 muldiv.scala 79:14]
  wire [63:0] _GEN_25 = _T_1 ? _GEN_17 : 64'h0; // @[Conditional.scala 39:67 muldiv.scala 77:12]
  wire [63:0] _GEN_26 = _T_1 ? _GEN_18 : 64'h0; // @[Conditional.scala 39:67 muldiv.scala 78:12]
  assign io_qua = _T ? 64'h0 : _GEN_25; // @[Conditional.scala 40:58 muldiv.scala 77:12]
  assign io_rem = _T ? 64'h0 : _GEN_26; // @[Conditional.scala 40:58 muldiv.scala 78:12]
  assign io_valid = _T ? 1'h0 : _GEN_24; // @[Conditional.scala 40:58 muldiv.scala 79:14]
  always @(posedge clock) begin
    if (reset) begin // @[muldiv.scala 67:27]
      quatient <= 64'h0; // @[muldiv.scala 67:27]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_en) begin // @[muldiv.scala 82:24]
        quatient <= 64'h0; // @[muldiv.scala 89:26]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (iter <= 7'h40) begin // @[muldiv.scala 94:39]
        quatient <= _GEN_8;
      end
    end
    if (reset) begin // @[muldiv.scala 68:26]
      val1 <= 128'h0; // @[muldiv.scala 68:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_en) begin // @[muldiv.scala 82:24]
        val1 <= _val1_T_6; // @[muldiv.scala 84:22]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (iter <= 7'h40) begin // @[muldiv.scala 94:39]
        val1 <= _GEN_9;
      end
    end
    if (reset) begin // @[muldiv.scala 69:26]
      val2 <= 128'h0; // @[muldiv.scala 69:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_en) begin // @[muldiv.scala 82:24]
        val2 <= _val2_T_6; // @[muldiv.scala 85:22]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (iter <= 7'h40) begin // @[muldiv.scala 94:39]
        val2 <= _GEN_10;
      end
    end
    if (reset) begin // @[muldiv.scala 70:27]
      qua_sign <= 1'h0; // @[muldiv.scala 70:27]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_en) begin // @[muldiv.scala 82:24]
        qua_sign <= io_sign & (io_a[63] != io_b[63] & io_b != 64'h0); // @[muldiv.scala 86:26]
      end
    end
    if (reset) begin // @[muldiv.scala 71:27]
      rem_sign <= 1'h0; // @[muldiv.scala 71:27]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_en) begin // @[muldiv.scala 82:24]
        rem_sign <= _val1_T_2; // @[muldiv.scala 87:26]
      end
    end
    if (reset) begin // @[muldiv.scala 72:26]
      iter <= 7'h0; // @[muldiv.scala 72:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_en) begin // @[muldiv.scala 82:24]
        iter <= 7'h0; // @[muldiv.scala 90:22]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (iter <= 7'h40) begin // @[muldiv.scala 94:39]
        iter <= _iter_T_1; // @[muldiv.scala 95:22]
      end
    end
    if (reset) begin // @[muldiv.scala 73:28]
      pre_alu64 <= 1'h0; // @[muldiv.scala 73:28]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_en) begin // @[muldiv.scala 82:24]
        pre_alu64 <= io_alu64; // @[muldiv.scala 88:27]
      end
    end
    if (reset) begin // @[muldiv.scala 75:24]
      state <= 2'h0; // @[muldiv.scala 75:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_en) begin // @[muldiv.scala 82:24]
        state <= 2'h1; // @[muldiv.scala 83:23]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (!(iter <= 7'h40)) begin // @[muldiv.scala 94:39]
        state <= 2'h0; // @[muldiv.scala 105:23]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  quatient = _RAND_0[63:0];
  _RAND_1 = {4{`RANDOM}};
  val1 = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  val2 = _RAND_2[127:0];
  _RAND_3 = {1{`RANDOM}};
  qua_sign = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  rem_sign = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  iter = _RAND_5[6:0];
  _RAND_6 = {1{`RANDOM}};
  pre_alu64 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_ALU(
  input         clock,
  input         reset,
  input  [4:0]  io_alu_op,
  input  [63:0] io_val1,
  input  [63:0] io_val2,
  input         io_alu64,
  input         io_en,
  output [63:0] io_out,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  multiplier_clock; // @[alu.scala 40:28]
  wire  multiplier_reset; // @[alu.scala 40:28]
  wire [63:0] multiplier_io_a; // @[alu.scala 40:28]
  wire [63:0] multiplier_io_b; // @[alu.scala 40:28]
  wire [4:0] multiplier_io_aluop; // @[alu.scala 40:28]
  wire  multiplier_io_en; // @[alu.scala 40:28]
  wire [63:0] multiplier_io_out; // @[alu.scala 40:28]
  wire  multiplier_io_valid; // @[alu.scala 40:28]
  wire  divider_clock; // @[alu.scala 41:28]
  wire  divider_reset; // @[alu.scala 41:28]
  wire  divider_io_alu64; // @[alu.scala 41:28]
  wire [63:0] divider_io_a; // @[alu.scala 41:28]
  wire [63:0] divider_io_b; // @[alu.scala 41:28]
  wire  divider_io_sign; // @[alu.scala 41:28]
  wire  divider_io_en; // @[alu.scala 41:28]
  wire [63:0] divider_io_qua; // @[alu.scala 41:28]
  wire [63:0] divider_io_rem; // @[alu.scala 41:28]
  wire  divider_io_valid; // @[alu.scala 41:28]
  reg [4:0] pre_aluop; // @[alu.scala 43:28]
  reg [1:0] state; // @[alu.scala 44:24]
  wire  _div_type_T_1 = 5'h11 == io_alu_op; // @[Lookup.scala 31:38]
  wire  _div_type_T_3 = 5'h12 == io_alu_op; // @[Lookup.scala 31:38]
  wire  _div_type_T_5 = 5'h13 == io_alu_op; // @[Lookup.scala 31:38]
  wire  _div_type_T_13 = _div_type_T_3 ? 1'h0 : _div_type_T_5; // @[Lookup.scala 33:37]
  wire  _T = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_7 = io_alu_op == 5'hd | io_alu_op == 5'he | io_alu_op == 5'hf | io_alu_op == 5'h10; // @[alu.scala 63:97]
  wire  _T_14 = io_alu_op == 5'h11 | io_alu_op == 5'h12 | io_alu_op == 5'h13 | io_alu_op == 5'h14; // @[alu.scala 66:102]
  wire [63:0] _alu_val_T_1 = io_val1 + io_val2; // @[alu.scala 75:49]
  wire [63:0] _alu_val_T_2 = io_val1 ^ io_val2; // @[alu.scala 76:49]
  wire [63:0] _alu_val_T_3 = io_val1 | io_val2; // @[alu.scala 77:49]
  wire [63:0] _alu_val_T_4 = io_val1 & io_val2; // @[alu.scala 78:49]
  wire [126:0] _GEN_33 = {{63'd0}, io_val1}; // @[alu.scala 79:49]
  wire [126:0] _alu_val_T_6 = _GEN_33 << io_val2[5:0]; // @[alu.scala 79:49]
  wire [63:0] _alu_val_T_8 = io_val1 >> io_val2[5:0]; // @[alu.scala 80:63]
  wire [31:0] _alu_val_T_11 = io_val1[31:0] >> io_val2[5:0]; // @[alu.scala 80:104]
  wire [63:0] _alu_val_T_12 = io_alu64 ? _alu_val_T_8 : {{32'd0}, _alu_val_T_11}; // @[alu.scala 80:43]
  wire [63:0] _alu_val_T_16 = $signed(io_val1) >>> io_val2[5:0]; // @[alu.scala 81:87]
  wire [31:0] _alu_val_T_18 = io_val1[31:0]; // @[alu.scala 81:112]
  wire [31:0] _alu_val_T_21 = $signed(_alu_val_T_18) >>> io_val2[5:0]; // @[alu.scala 81:136]
  wire [63:0] _alu_val_T_22 = io_alu64 ? _alu_val_T_16 : {{32'd0}, _alu_val_T_21}; // @[alu.scala 81:43]
  wire [63:0] _alu_val_T_24 = io_val1 - io_val2; // @[alu.scala 82:49]
  wire  _alu_val_T_27 = $signed(io_val1) < $signed(io_val2); // @[alu.scala 83:59]
  wire  _alu_val_T_29 = io_val1 < io_val2; // @[alu.scala 84:52]
  wire [63:0] _alu_val_T_31 = ~io_val1; // @[alu.scala 85:42]
  wire [63:0] _alu_val_T_32 = _alu_val_T_31 & io_val2; // @[alu.scala 85:52]
  wire [63:0] _alu_val_T_36 = 5'h1 == io_alu_op ? io_val1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _alu_val_T_38 = 5'h2 == io_alu_op ? io_val2 : _alu_val_T_36; // @[Mux.scala 80:57]
  wire [63:0] _alu_val_T_40 = 5'h3 == io_alu_op ? _alu_val_T_1 : _alu_val_T_38; // @[Mux.scala 80:57]
  wire [63:0] _alu_val_T_42 = 5'h4 == io_alu_op ? _alu_val_T_2 : _alu_val_T_40; // @[Mux.scala 80:57]
  wire [63:0] _alu_val_T_44 = 5'h5 == io_alu_op ? _alu_val_T_3 : _alu_val_T_42; // @[Mux.scala 80:57]
  wire [63:0] _alu_val_T_46 = 5'h6 == io_alu_op ? _alu_val_T_4 : _alu_val_T_44; // @[Mux.scala 80:57]
  wire [126:0] _alu_val_T_48 = 5'h7 == io_alu_op ? _alu_val_T_6 : {{63'd0}, _alu_val_T_46}; // @[Mux.scala 80:57]
  wire [126:0] _alu_val_T_50 = 5'h8 == io_alu_op ? {{63'd0}, _alu_val_T_12} : _alu_val_T_48; // @[Mux.scala 80:57]
  wire [126:0] _alu_val_T_52 = 5'h9 == io_alu_op ? {{63'd0}, _alu_val_T_22} : _alu_val_T_50; // @[Mux.scala 80:57]
  wire [126:0] _alu_val_T_54 = 5'ha == io_alu_op ? {{63'd0}, _alu_val_T_24} : _alu_val_T_52; // @[Mux.scala 80:57]
  wire [126:0] _alu_val_T_56 = 5'hb == io_alu_op ? {{126'd0}, _alu_val_T_27} : _alu_val_T_54; // @[Mux.scala 80:57]
  wire [126:0] _alu_val_T_58 = 5'hc == io_alu_op ? {{126'd0}, _alu_val_T_29} : _alu_val_T_56; // @[Mux.scala 80:57]
  wire [126:0] alu_val = 5'h15 == io_alu_op ? {{63'd0}, _alu_val_T_32} : _alu_val_T_58; // @[Mux.scala 80:57]
  wire [1:0] _GEN_1 = io_alu_op == 5'h11 | io_alu_op == 5'h12 | io_alu_op == 5'h13 | io_alu_op == 5'h14 ? 2'h2 : state; // @[alu.scala 66:129 alu.scala 68:27 alu.scala 44:24]
  wire [126:0] _GEN_2 = io_alu_op == 5'h11 | io_alu_op == 5'h12 | io_alu_op == 5'h13 | io_alu_op == 5'h14 ? 127'h0 :
    alu_val; // @[alu.scala 66:129 alu.scala 57:14 alu.scala 87:28]
  wire  _GEN_3 = io_alu_op == 5'h11 | io_alu_op == 5'h12 | io_alu_op == 5'h13 | io_alu_op == 5'h14 ? 1'h0 : 1'h1; // @[alu.scala 66:129 alu.scala 56:14 alu.scala 88:30]
  wire  _GEN_6 = io_alu_op == 5'hd | io_alu_op == 5'he | io_alu_op == 5'hf | io_alu_op == 5'h10 ? 1'h0 : _T_14; // @[alu.scala 63:125 alu.scala 55:25]
  wire [126:0] _GEN_7 = io_alu_op == 5'hd | io_alu_op == 5'he | io_alu_op == 5'hf | io_alu_op == 5'h10 ? 127'h0 : _GEN_2
    ; // @[alu.scala 63:125 alu.scala 57:14]
  wire  _GEN_8 = io_alu_op == 5'hd | io_alu_op == 5'he | io_alu_op == 5'hf | io_alu_op == 5'h10 ? 1'h0 : _GEN_3; // @[alu.scala 63:125 alu.scala 56:14]
  wire  _GEN_10 = io_en & _T_7; // @[alu.scala 61:24 alu.scala 48:25]
  wire  _GEN_12 = io_en & _GEN_6; // @[alu.scala 61:24 alu.scala 55:25]
  wire [126:0] _GEN_13 = io_en ? _GEN_7 : 127'h0; // @[alu.scala 61:24 alu.scala 57:14]
  wire  _GEN_14 = io_en & _GEN_8; // @[alu.scala 61:24 alu.scala 56:14]
  wire  _T_15 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire [63:0] _GEN_15 = multiplier_io_valid ? multiplier_io_out : 64'h0; // @[alu.scala 93:38 alu.scala 94:24 alu.scala 57:14]
  wire  _GEN_16 = multiplier_io_valid; // @[alu.scala 93:38 alu.scala 95:26 alu.scala 56:14]
  wire  _T_16 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [63:0] _io_out_T_3 = pre_aluop == 5'h11 | pre_aluop == 5'h12 ? divider_io_qua : divider_io_rem; // @[alu.scala 101:30]
  wire [63:0] _GEN_18 = divider_io_valid ? _io_out_T_3 : 64'h0; // @[alu.scala 100:35 alu.scala 101:24 alu.scala 57:14]
  wire  _GEN_19 = divider_io_valid; // @[alu.scala 100:35 alu.scala 102:26 alu.scala 56:14]
  wire [1:0] _GEN_20 = divider_io_valid ? 2'h0 : state; // @[alu.scala 100:35 alu.scala 103:23 alu.scala 44:24]
  wire [63:0] _GEN_21 = _T_16 ? _GEN_18 : 64'h0; // @[Conditional.scala 39:67 alu.scala 57:14]
  wire  _GEN_22 = _T_16 & _GEN_19; // @[Conditional.scala 39:67 alu.scala 56:14]
  wire [63:0] _GEN_24 = _T_15 ? _GEN_15 : _GEN_21; // @[Conditional.scala 39:67]
  wire  _GEN_25 = _T_15 ? _GEN_16 : _GEN_22; // @[Conditional.scala 39:67]
  wire [126:0] _GEN_31 = _T ? _GEN_13 : {{63'd0}, _GEN_24}; // @[Conditional.scala 40:58]
  ysyx_210539_MUL multiplier ( // @[alu.scala 40:28]
    .clock(multiplier_clock),
    .reset(multiplier_reset),
    .io_a(multiplier_io_a),
    .io_b(multiplier_io_b),
    .io_aluop(multiplier_io_aluop),
    .io_en(multiplier_io_en),
    .io_out(multiplier_io_out),
    .io_valid(multiplier_io_valid)
  );
  ysyx_210539_DIV divider ( // @[alu.scala 41:28]
    .clock(divider_clock),
    .reset(divider_reset),
    .io_alu64(divider_io_alu64),
    .io_a(divider_io_a),
    .io_b(divider_io_b),
    .io_sign(divider_io_sign),
    .io_en(divider_io_en),
    .io_qua(divider_io_qua),
    .io_rem(divider_io_rem),
    .io_valid(divider_io_valid)
  );
  assign io_out = _GEN_31[63:0];
  assign io_valid = _T ? _GEN_14 : _GEN_25; // @[Conditional.scala 40:58]
  assign multiplier_clock = clock;
  assign multiplier_reset = reset;
  assign multiplier_io_a = io_val1; // @[alu.scala 46:25]
  assign multiplier_io_b = io_val2; // @[alu.scala 47:25]
  assign multiplier_io_aluop = io_alu_op; // @[alu.scala 49:26]
  assign multiplier_io_en = _T & _GEN_10; // @[Conditional.scala 40:58 alu.scala 48:25]
  assign divider_clock = clock;
  assign divider_reset = reset;
  assign divider_io_alu64 = io_alu64; // @[alu.scala 51:25]
  assign divider_io_a = io_val1; // @[alu.scala 52:25]
  assign divider_io_b = io_val2; // @[alu.scala 53:25]
  assign divider_io_sign = _div_type_T_1 | _div_type_T_13; // @[Lookup.scala 33:37]
  assign divider_io_en = _T & _GEN_12; // @[Conditional.scala 40:58 alu.scala 55:25]
  always @(posedge clock) begin
    if (reset) begin // @[alu.scala 43:28]
      pre_aluop <= 5'h0; // @[alu.scala 43:28]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_en) begin // @[alu.scala 61:24]
        pre_aluop <= io_alu_op; // @[alu.scala 62:27]
      end
    end
    if (reset) begin // @[alu.scala 44:24]
      state <= 2'h0; // @[alu.scala 44:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_en) begin // @[alu.scala 61:24]
        if (io_alu_op == 5'hd | io_alu_op == 5'he | io_alu_op == 5'hf | io_alu_op == 5'h10) begin // @[alu.scala 63:125]
          state <= 2'h1; // @[alu.scala 65:27]
        end else begin
          state <= _GEN_1;
        end
      end
    end else if (_T_15) begin // @[Conditional.scala 39:67]
      if (multiplier_io_valid) begin // @[alu.scala 93:38]
        state <= 2'h0; // @[alu.scala 96:23]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_20;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pre_aluop = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_BranchALU(
  input  [63:0] io_val1,
  input  [63:0] io_val2,
  input  [2:0]  io_brType,
  output        io_is_jmp
);
  wire  _io_is_jmp_T = io_val1 == io_val2; // @[alu.scala 119:29]
  wire  _io_is_jmp_T_1 = io_val1 != io_val2; // @[alu.scala 120:29]
  wire  _io_is_jmp_T_4 = $signed(io_val1) < $signed(io_val2); // @[alu.scala 121:36]
  wire  _io_is_jmp_T_7 = $signed(io_val1) >= $signed(io_val2); // @[alu.scala 122:36]
  wire  _io_is_jmp_T_8 = io_val1 < io_val2; // @[alu.scala 123:29]
  wire  _io_is_jmp_T_9 = io_val1 >= io_val2; // @[alu.scala 124:29]
  wire  _io_is_jmp_T_13 = 3'h1 == io_brType ? _io_is_jmp_T_1 : 3'h0 == io_brType & _io_is_jmp_T; // @[Mux.scala 80:57]
  wire  _io_is_jmp_T_15 = 3'h4 == io_brType ? _io_is_jmp_T_4 : _io_is_jmp_T_13; // @[Mux.scala 80:57]
  wire  _io_is_jmp_T_17 = 3'h5 == io_brType ? _io_is_jmp_T_7 : _io_is_jmp_T_15; // @[Mux.scala 80:57]
  wire  _io_is_jmp_T_19 = 3'h6 == io_brType ? _io_is_jmp_T_8 : _io_is_jmp_T_17; // @[Mux.scala 80:57]
  assign io_is_jmp = 3'h7 == io_brType ? _io_is_jmp_T_9 : _io_is_jmp_T_19; // @[Mux.scala 80:57]
endmodule
module ysyx_210539_Execute(
  input         clock,
  input         reset,
  input  [31:0] io_rr2ex_inst,
  input  [63:0] io_rr2ex_pc,
  input  [63:0] io_rr2ex_excep_cause,
  input  [63:0] io_rr2ex_excep_tval,
  input         io_rr2ex_excep_en,
  input  [63:0] io_rr2ex_excep_pc,
  input  [1:0]  io_rr2ex_excep_etype,
  input  [4:0]  io_rr2ex_ctrl_aluOp,
  input         io_rr2ex_ctrl_aluWidth,
  input  [4:0]  io_rr2ex_ctrl_dcMode,
  input         io_rr2ex_ctrl_writeRegEn,
  input         io_rr2ex_ctrl_writeCSREn,
  input  [2:0]  io_rr2ex_ctrl_brType,
  input  [63:0] io_rr2ex_rs1_d,
  input  [11:0] io_rr2ex_rs2,
  input  [63:0] io_rr2ex_rs2_d,
  input  [4:0]  io_rr2ex_dst,
  input  [63:0] io_rr2ex_dst_d,
  input  [11:0] io_rr2ex_rcsr_id,
  input  [1:0]  io_rr2ex_jmp_type,
  input  [1:0]  io_rr2ex_special,
  input  [1:0]  io_rr2ex_indi,
  output        io_rr2ex_drop,
  output        io_rr2ex_stall,
  input         io_rr2ex_recov,
  input         io_rr2ex_valid,
  output        io_rr2ex_ready,
  output [31:0] io_ex2mem_inst,
  output [63:0] io_ex2mem_pc,
  output [63:0] io_ex2mem_excep_cause,
  output [63:0] io_ex2mem_excep_tval,
  output        io_ex2mem_excep_en,
  output [63:0] io_ex2mem_excep_pc,
  output [1:0]  io_ex2mem_excep_etype,
  output [4:0]  io_ex2mem_ctrl_dcMode,
  output        io_ex2mem_ctrl_writeRegEn,
  output        io_ex2mem_ctrl_writeCSREn,
  output [63:0] io_ex2mem_mem_addr,
  output [63:0] io_ex2mem_mem_data,
  output [11:0] io_ex2mem_csr_id,
  output [63:0] io_ex2mem_csr_d,
  output [4:0]  io_ex2mem_dst,
  output [63:0] io_ex2mem_dst_d,
  output [11:0] io_ex2mem_rcsr_id,
  output [1:0]  io_ex2mem_special,
  output [1:0]  io_ex2mem_indi,
  input         io_ex2mem_drop,
  input         io_ex2mem_stall,
  output        io_ex2mem_recov,
  output        io_ex2mem_valid,
  input         io_ex2mem_ready,
  output [4:0]  io_d_ex_id,
  output [63:0] io_d_ex_data,
  output [1:0]  io_d_ex_state,
  output [63:0] io_ex2if_seq_pc,
  output        io_ex2if_valid,
  input  [63:0] io_updateNextPc_seq_pc,
  input         io_updateNextPc_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  wire  alu_clock; // @[execute.scala 27:25]
  wire  alu_reset; // @[execute.scala 27:25]
  wire [4:0] alu_io_alu_op; // @[execute.scala 27:25]
  wire [63:0] alu_io_val1; // @[execute.scala 27:25]
  wire [63:0] alu_io_val2; // @[execute.scala 27:25]
  wire  alu_io_alu64; // @[execute.scala 27:25]
  wire  alu_io_en; // @[execute.scala 27:25]
  wire [63:0] alu_io_out; // @[execute.scala 27:25]
  wire  alu_io_valid; // @[execute.scala 27:25]
  wire [63:0] branchAlu_io_val1; // @[execute.scala 153:27]
  wire [63:0] branchAlu_io_val2; // @[execute.scala 153:27]
  wire [2:0] branchAlu_io_brType; // @[execute.scala 153:27]
  wire  branchAlu_io_is_jmp; // @[execute.scala 153:27]
  reg  drop_r; // @[execute.scala 21:25]
  reg  stall_r; // @[execute.scala 22:26]
  wire  drop_in = drop_r | io_ex2mem_drop; // @[execute.scala 24:26]
  wire  _io_rr2ex_stall_T = ~io_ex2mem_drop; // @[execute.scala 26:55]
  reg [31:0] inst_r; // @[execute.scala 28:30]
  reg [63:0] pc_r; // @[execute.scala 29:30]
  reg [63:0] excep_r_cause; // @[execute.scala 30:30]
  reg [63:0] excep_r_tval; // @[execute.scala 30:30]
  reg  excep_r_en; // @[execute.scala 30:30]
  reg [63:0] excep_r_pc; // @[execute.scala 30:30]
  reg [1:0] excep_r_etype; // @[execute.scala 30:30]
  reg [4:0] ctrl_r_dcMode; // @[execute.scala 31:30]
  reg  ctrl_r_writeRegEn; // @[execute.scala 31:30]
  reg  ctrl_r_writeCSREn; // @[execute.scala 31:30]
  reg [63:0] mem_addr_r; // @[execute.scala 32:30]
  reg [63:0] mem_data_r; // @[execute.scala 33:30]
  reg [11:0] csr_id_r; // @[execute.scala 34:30]
  reg [63:0] csr_d_r; // @[execute.scala 35:30]
  reg [4:0] dst_r; // @[execute.scala 36:30]
  reg [63:0] dst_d_r; // @[execute.scala 37:30]
  reg [11:0] rcsr_id_r; // @[execute.scala 38:30]
  reg [1:0] special_r; // @[execute.scala 39:30]
  reg  alu64_r; // @[execute.scala 40:30]
  reg [1:0] indi_r; // @[execute.scala 41:30]
  reg [63:0] next_pc_r; // @[execute.scala 42:30]
  reg  recov_r; // @[execute.scala 43:30]
  reg  valid_r; // @[execute.scala 44:30]
  wire  hs_in = io_rr2ex_ready & io_rr2ex_valid; // @[execute.scala 46:34]
  wire  hs_out = io_ex2mem_ready & io_ex2mem_valid; // @[execute.scala 47:35]
  wire  alu64 = ~io_rr2ex_ctrl_aluWidth; // @[execute.scala 48:40]
  wire  _signed_dr_T = ~alu64; // @[execute.scala 51:23]
  wire  signed_dr = ~alu64 & (io_rr2ex_ctrl_aluOp == 5'h11 | io_rr2ex_ctrl_aluOp == 5'h13); // @[execute.scala 51:30]
  wire  unsigned_dr = _signed_dr_T & (io_rr2ex_ctrl_aluOp == 5'h12 | io_rr2ex_ctrl_aluOp == 5'h14); // @[execute.scala 52:30]
  wire [31:0] val1_lo = io_rr2ex_rs1_d[31:0]; // @[common.scala 712:29]
  wire [63:0] _val1_T = {32'h0,val1_lo}; // @[Cat.scala 30:58]
  wire [31:0] val1_hi = io_rr2ex_rs1_d[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _val1_T_3 = {val1_hi,val1_lo}; // @[Cat.scala 30:58]
  wire [63:0] _val1_T_4 = signed_dr ? _val1_T_3 : io_rr2ex_rs1_d; // @[Mux.scala 47:69]
  wire  is_shift = io_rr2ex_ctrl_aluOp == 5'h7 | io_rr2ex_ctrl_aluOp == 5'h8 | io_rr2ex_ctrl_aluOp == 5'h9; // @[execute.scala 58:59]
  wire [31:0] val2_lo = io_rr2ex_rs2_d[31:0]; // @[common.scala 712:29]
  wire [63:0] _val2_T = {32'h0,val2_lo}; // @[Cat.scala 30:58]
  wire [31:0] val2_hi = io_rr2ex_rs2_d[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _val2_T_3 = {val2_hi,val2_lo}; // @[Cat.scala 30:58]
  wire [4:0] val2_lo_2 = io_rr2ex_rs2_d[4:0]; // @[execute.scala 62:85]
  wire [5:0] _val2_T_5 = {1'h0,val2_lo_2}; // @[Cat.scala 30:58]
  wire [5:0] _val2_T_6 = alu64 ? io_rr2ex_rs2_d[5:0] : _val2_T_5; // @[execute.scala 62:28]
  wire [63:0] _val2_T_7 = is_shift ? {{58'd0}, _val2_T_6} : io_rr2ex_rs2_d; // @[Mux.scala 47:69]
  wire [63:0] _val2_T_8 = signed_dr ? _val2_T_3 : _val2_T_7; // @[Mux.scala 47:69]
  wire  cur_alu64 = hs_in ? alu64 : alu64_r; // @[execute.scala 70:26]
  wire [63:0] _alu_out_T = alu_io_out; // @[execute.scala 71:44]
  wire [31:0] alu_out_hi = alu_io_out[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] alu_out_lo = alu_io_out[31:0]; // @[common.scala 709:40]
  wire [63:0] _alu_out_T_3 = {alu_out_hi,alu_out_lo}; // @[Cat.scala 30:58]
  wire [63:0] alu_out = cur_alu64 ? _alu_out_T : _alu_out_T_3; // @[execute.scala 71:22]
  wire [63:0] _wdata_T_1 = io_rr2ex_ctrl_writeCSREn ? io_rr2ex_rs2_d : alu_out; // @[Mux.scala 47:69]
  wire [63:0] wdata = io_rr2ex_ctrl_dcMode[3] ? io_rr2ex_dst_d : _wdata_T_1; // @[Mux.scala 47:69]
  wire [63:0] _memAlign_ans_T = alu_out & 64'h1; // @[common.scala 329:27]
  wire  _memAlign_ans_T_1 = _memAlign_ans_T == 64'h0; // @[common.scala 329:36]
  wire [63:0] _memAlign_ans_T_2 = alu_out & 64'h3; // @[common.scala 330:27]
  wire  _memAlign_ans_T_3 = _memAlign_ans_T_2 == 64'h0; // @[common.scala 330:36]
  wire [63:0] _memAlign_ans_T_4 = alu_out & 64'h7; // @[common.scala 331:27]
  wire  _memAlign_ans_T_5 = _memAlign_ans_T_4 == 64'h0; // @[common.scala 331:36]
  wire  _memAlign_ans_T_7 = 2'h1 == io_rr2ex_ctrl_dcMode[1:0] ? _memAlign_ans_T_1 : 1'h1; // @[Mux.scala 80:57]
  wire  _memAlign_ans_T_9 = 2'h2 == io_rr2ex_ctrl_dcMode[1:0] ? _memAlign_ans_T_3 : _memAlign_ans_T_7; // @[Mux.scala 80:57]
  wire  memAlign_ans = 2'h3 == io_rr2ex_ctrl_dcMode[1:0] ? _memAlign_ans_T_5 : _memAlign_ans_T_9; // @[Mux.scala 80:57]
  wire  memAlign = io_rr2ex_ctrl_dcMode == 5'h0 | memAlign_ans; // @[execute.scala 85:54]
  wire  _T_1 = ~memAlign; // @[execute.scala 105:14]
  wire [2:0] _excep_r_cause_T_1 = io_rr2ex_ctrl_dcMode[3] ? 3'h6 : 3'h4; // @[execute.scala 108:33]
  wire  _GEN_11 = ~memAlign | io_rr2ex_excep_en; // @[execute.scala 105:24 execute.scala 110:25 execute.scala 89:21]
  wire  _GEN_15 = ~memAlign | io_rr2ex_recov; // @[execute.scala 105:24 execute.scala 83:54 execute.scala 101:21]
  wire [63:0] _GEN_34 = hs_in ? wdata : dst_d_r; // @[execute.scala 86:16 execute.scala 96:21 execute.scala 37:30]
  wire  _GEN_40 = hs_in & _T_1; // @[execute.scala 86:16 execute.scala 23:12]
  reg  state; // @[execute.scala 118:24]
  reg  drop_alu; // @[execute.scala 119:27]
  wire  _T_2 = ~drop_in; // @[execute.scala 120:10]
  wire  _GEN_42 = (valid_r | state) & ~hs_out ? 1'h0 : io_rr2ex_valid; // @[execute.scala 121:54 execute.scala 116:21]
  wire  _GEN_44 = hs_out ? 1'h0 : valid_r; // @[execute.scala 134:31 execute.scala 135:25 execute.scala 44:30]
  wire  _GEN_45 = hs_in | _GEN_44; // @[execute.scala 132:30 execute.scala 133:25]
  wire  _GEN_46 = hs_in & ~alu_io_valid ? 1'h0 : _GEN_45; // @[execute.scala 129:41 execute.scala 130:25]
  wire  _GEN_47 = hs_in & ~alu_io_valid | state; // @[execute.scala 129:41 execute.scala 131:23 execute.scala 118:24]
  wire  _GEN_48 = ~state ? _GEN_46 : valid_r; // @[execute.scala 128:30 execute.scala 44:30]
  wire  _GEN_49 = ~state ? _GEN_47 : state; // @[execute.scala 128:30 execute.scala 118:24]
  wire  _GEN_52 = alu_io_valid ? ~drop_alu : _GEN_48; // @[execute.scala 139:31 execute.scala 142:29]
  wire  _GEN_56 = state ? _GEN_52 : _GEN_48; // @[execute.scala 138:33]
  wire  _GEN_58 = state | drop_alu; // @[execute.scala 148:30 execute.scala 149:22 execute.scala 119:27]
  wire  _GEN_59 = _io_rr2ex_stall_T & _GEN_56; // @[execute.scala 127:26 execute.scala 147:17]
  reg [63:0] forceJmp_seq_pc; // @[execute.scala 154:27]
  reg  forceJmp_valid; // @[execute.scala 154:27]
  wire  real_is_target = 2'h2 == io_rr2ex_jmp_type ? branchAlu_io_is_jmp : 2'h1 == io_rr2ex_jmp_type; // @[Mux.scala 80:57]
  wire  _real_target_T = io_rr2ex_jmp_type == 2'h3; // @[execute.scala 164:28]
  wire  _real_target_T_1 = ~real_is_target; // @[execute.scala 165:10]
  wire [2:0] _real_target_T_4 = io_rr2ex_inst[1:0] == 2'h3 ? 3'h4 : 3'h2; // @[execute.scala 165:62]
  wire [63:0] _GEN_72 = {{61'd0}, _real_target_T_4}; // @[execute.scala 165:57]
  wire [63:0] _real_target_T_6 = io_rr2ex_pc + _GEN_72; // @[execute.scala 165:57]
  wire  _real_target_T_7 = io_rr2ex_jmp_type == 2'h1; // @[execute.scala 166:28]
  wire [63:0] _real_target_T_9 = io_rr2ex_rs1_d + io_rr2ex_dst_d; // @[execute.scala 166:60]
  wire [63:0] _real_target_T_10 = _real_target_T_7 ? _real_target_T_9 : io_rr2ex_dst_d; // @[Mux.scala 47:69]
  wire [63:0] _real_target_T_11 = _real_target_T_1 ? _real_target_T_6 : _real_target_T_10; // @[Mux.scala 47:69]
  wire  _T_18 = hs_in & ~io_rr2ex_excep_en & real_is_target & io_rr2ex_jmp_type != 2'h0; // @[execute.scala 174:60]
  wire  _GEN_66 = hs_in & ~io_rr2ex_excep_en & real_is_target & io_rr2ex_jmp_type != 2'h0 | _GEN_40; // @[execute.scala 174:92 execute.scala 177:21]
  wire  _GEN_68 = _T_2 & _T_18; // @[execute.scala 173:19 execute.scala 155:20]
  wire [1:0] _io_d_ex_state_T_3 = ctrl_r_writeRegEn ? 2'h1 : 2'h0; // @[execute.scala 189:91]
  wire [1:0] _io_d_ex_state_T_4 = ctrl_r_dcMode[2] | indi_r[1] ? 2'h2 : _io_d_ex_state_T_3; // @[execute.scala 189:31]
  wire [1:0] _GEN_70 = state ? 2'h2 : 2'h0; // @[execute.scala 190:32 execute.scala 191:25 execute.scala 187:20]
  ysyx_210539_ALU alu ( // @[execute.scala 27:25]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_alu_op(alu_io_alu_op),
    .io_val1(alu_io_val1),
    .io_val2(alu_io_val2),
    .io_alu64(alu_io_alu64),
    .io_en(alu_io_en),
    .io_out(alu_io_out),
    .io_valid(alu_io_valid)
  );
  ysyx_210539_BranchALU branchAlu ( // @[execute.scala 153:27]
    .io_val1(branchAlu_io_val1),
    .io_val2(branchAlu_io_val2),
    .io_brType(branchAlu_io_brType),
    .io_is_jmp(branchAlu_io_is_jmp)
  );
  assign io_rr2ex_drop = drop_r | io_ex2mem_drop; // @[execute.scala 24:26]
  assign io_rr2ex_stall = io_ex2mem_stall | stall_r & ~io_ex2mem_drop; // @[execute.scala 26:40]
  assign io_rr2ex_ready = ~drop_in & _GEN_42; // @[execute.scala 120:19 execute.scala 116:21]
  assign io_ex2mem_inst = inst_r; // @[execute.scala 195:25]
  assign io_ex2mem_pc = pc_r; // @[execute.scala 196:25]
  assign io_ex2mem_excep_cause = excep_r_cause; // @[execute.scala 197:25]
  assign io_ex2mem_excep_tval = excep_r_tval; // @[execute.scala 197:25]
  assign io_ex2mem_excep_en = excep_r_en; // @[execute.scala 197:25]
  assign io_ex2mem_excep_pc = excep_r_pc; // @[execute.scala 197:25]
  assign io_ex2mem_excep_etype = excep_r_etype; // @[execute.scala 197:25]
  assign io_ex2mem_ctrl_dcMode = ctrl_r_dcMode; // @[execute.scala 198:25]
  assign io_ex2mem_ctrl_writeRegEn = ctrl_r_writeRegEn; // @[execute.scala 198:25]
  assign io_ex2mem_ctrl_writeCSREn = ctrl_r_writeCSREn; // @[execute.scala 198:25]
  assign io_ex2mem_mem_addr = mem_addr_r; // @[execute.scala 199:25]
  assign io_ex2mem_mem_data = mem_data_r; // @[execute.scala 200:25]
  assign io_ex2mem_csr_id = csr_id_r; // @[execute.scala 201:25]
  assign io_ex2mem_csr_d = csr_d_r; // @[execute.scala 202:25]
  assign io_ex2mem_dst = dst_r; // @[execute.scala 203:25]
  assign io_ex2mem_dst_d = dst_d_r; // @[execute.scala 204:25]
  assign io_ex2mem_rcsr_id = rcsr_id_r; // @[execute.scala 205:25]
  assign io_ex2mem_special = special_r; // @[execute.scala 206:25]
  assign io_ex2mem_indi = indi_r; // @[execute.scala 207:25]
  assign io_ex2mem_recov = recov_r; // @[execute.scala 209:25]
  assign io_ex2mem_valid = valid_r; // @[execute.scala 208:25]
  assign io_d_ex_id = dst_r; // @[execute.scala 185:20]
  assign io_d_ex_data = dst_d_r; // @[execute.scala 186:20]
  assign io_d_ex_state = valid_r ? _io_d_ex_state_T_4 : _GEN_70; // @[execute.scala 188:18 execute.scala 189:25]
  assign io_ex2if_seq_pc = forceJmp_seq_pc; // @[execute.scala 180:21]
  assign io_ex2if_valid = forceJmp_valid & _io_rr2ex_stall_T; // @[execute.scala 181:39]
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_alu_op = io_rr2ex_ctrl_aluOp; // @[execute.scala 65:21]
  assign alu_io_val1 = unsigned_dr ? _val1_T : _val1_T_4; // @[Mux.scala 47:69]
  assign alu_io_val2 = unsigned_dr ? _val2_T : _val2_T_8; // @[Mux.scala 47:69]
  assign alu_io_alu64 = ~io_rr2ex_ctrl_aluWidth; // @[execute.scala 48:40]
  assign alu_io_en = ~drop_in & _GEN_42; // @[execute.scala 120:19 execute.scala 116:21]
  assign branchAlu_io_val1 = unsigned_dr ? _val1_T : _val1_T_4; // @[Mux.scala 47:69]
  assign branchAlu_io_val2 = unsigned_dr ? _val2_T : _val2_T_8; // @[Mux.scala 47:69]
  assign branchAlu_io_brType = io_rr2ex_ctrl_brType; // @[execute.scala 158:25]
  always @(posedge clock) begin
    if (reset) begin // @[execute.scala 21:25]
      drop_r <= 1'h0; // @[execute.scala 21:25]
    end else if (_T_2) begin // @[execute.scala 173:19]
      drop_r <= _GEN_66;
    end else begin
      drop_r <= _GEN_40;
    end
    if (reset) begin // @[execute.scala 22:26]
      stall_r <= 1'h0; // @[execute.scala 22:26]
    end else begin
      stall_r <= _GEN_40;
    end
    if (reset) begin // @[execute.scala 28:30]
      inst_r <= 32'h0; // @[execute.scala 28:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      inst_r <= io_rr2ex_inst; // @[execute.scala 87:21]
    end
    if (reset) begin // @[execute.scala 29:30]
      pc_r <= 64'h0; // @[execute.scala 29:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      pc_r <= io_rr2ex_pc; // @[execute.scala 88:21]
    end
    if (reset) begin // @[execute.scala 30:30]
      excep_r_cause <= 64'h0; // @[execute.scala 30:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      if (~memAlign) begin // @[execute.scala 105:24]
        excep_r_cause <= {{61'd0}, _excep_r_cause_T_1}; // @[execute.scala 108:27]
      end else begin
        excep_r_cause <= io_rr2ex_excep_cause; // @[execute.scala 89:21]
      end
    end
    if (reset) begin // @[execute.scala 30:30]
      excep_r_tval <= 64'h0; // @[execute.scala 30:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      if (~memAlign) begin // @[execute.scala 105:24]
        if (cur_alu64) begin // @[execute.scala 71:22]
          excep_r_tval <= _alu_out_T;
        end else begin
          excep_r_tval <= _alu_out_T_3;
        end
      end else begin
        excep_r_tval <= io_rr2ex_excep_tval; // @[execute.scala 89:21]
      end
    end
    if (reset) begin // @[execute.scala 30:30]
      excep_r_en <= 1'h0; // @[execute.scala 30:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      excep_r_en <= _GEN_11;
    end
    if (reset) begin // @[execute.scala 30:30]
      excep_r_pc <= 64'h0; // @[execute.scala 30:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      if (~memAlign) begin // @[execute.scala 105:24]
        excep_r_pc <= io_rr2ex_pc; // @[execute.scala 111:25]
      end else if (io_rr2ex_excep_cause[63]) begin // @[execute.scala 102:39]
        excep_r_pc <= next_pc_r; // @[execute.scala 103:24]
      end else begin
        excep_r_pc <= io_rr2ex_excep_pc; // @[execute.scala 89:21]
      end
    end
    if (reset) begin // @[execute.scala 30:30]
      excep_r_etype <= 2'h0; // @[execute.scala 30:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      if (~memAlign) begin // @[execute.scala 105:24]
        excep_r_etype <= 2'h0; // @[execute.scala 112:27]
      end else begin
        excep_r_etype <= io_rr2ex_excep_etype; // @[execute.scala 89:21]
      end
    end
    if (reset) begin // @[execute.scala 31:30]
      ctrl_r_dcMode <= 5'h0; // @[execute.scala 31:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      if (~memAlign) begin // @[execute.scala 105:24]
        ctrl_r_dcMode <= 5'h0; // @[execute.scala 106:20]
      end else begin
        ctrl_r_dcMode <= io_rr2ex_ctrl_dcMode; // @[execute.scala 90:21]
      end
    end
    if (reset) begin // @[execute.scala 31:30]
      ctrl_r_writeRegEn <= 1'h0; // @[execute.scala 31:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      if (~memAlign) begin // @[execute.scala 105:24]
        ctrl_r_writeRegEn <= 1'h0; // @[execute.scala 106:20]
      end else begin
        ctrl_r_writeRegEn <= io_rr2ex_ctrl_writeRegEn; // @[execute.scala 90:21]
      end
    end
    if (reset) begin // @[execute.scala 31:30]
      ctrl_r_writeCSREn <= 1'h0; // @[execute.scala 31:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      if (~memAlign) begin // @[execute.scala 105:24]
        ctrl_r_writeCSREn <= 1'h0; // @[execute.scala 106:20]
      end else begin
        ctrl_r_writeCSREn <= io_rr2ex_ctrl_writeCSREn; // @[execute.scala 90:21]
      end
    end
    if (reset) begin // @[execute.scala 32:30]
      mem_addr_r <= 64'h0; // @[execute.scala 32:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      if (cur_alu64) begin // @[execute.scala 71:22]
        mem_addr_r <= _alu_out_T;
      end else begin
        mem_addr_r <= _alu_out_T_3;
      end
    end
    if (reset) begin // @[execute.scala 33:30]
      mem_data_r <= 64'h0; // @[execute.scala 33:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      if (io_rr2ex_ctrl_dcMode[3]) begin // @[Mux.scala 47:69]
        mem_data_r <= io_rr2ex_dst_d;
      end else if (io_rr2ex_ctrl_writeCSREn) begin // @[Mux.scala 47:69]
        mem_data_r <= io_rr2ex_rs2_d;
      end else begin
        mem_data_r <= alu_out;
      end
    end
    if (reset) begin // @[execute.scala 34:30]
      csr_id_r <= 12'h0; // @[execute.scala 34:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      csr_id_r <= io_rr2ex_rs2; // @[execute.scala 93:21]
    end
    if (reset) begin // @[execute.scala 35:30]
      csr_d_r <= 64'h0; // @[execute.scala 35:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      if (cur_alu64) begin // @[execute.scala 71:22]
        csr_d_r <= _alu_out_T;
      end else begin
        csr_d_r <= _alu_out_T_3;
      end
    end
    if (reset) begin // @[execute.scala 36:30]
      dst_r <= 5'h0; // @[execute.scala 36:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      dst_r <= io_rr2ex_dst; // @[execute.scala 95:21]
    end
    if (reset) begin // @[execute.scala 37:30]
      dst_d_r <= 64'h0; // @[execute.scala 37:30]
    end else if (_io_rr2ex_stall_T) begin // @[execute.scala 127:26]
      if (state) begin // @[execute.scala 138:33]
        if (alu_io_valid) begin // @[execute.scala 139:31]
          dst_d_r <= alu_out; // @[execute.scala 141:29]
        end else begin
          dst_d_r <= _GEN_34;
        end
      end else begin
        dst_d_r <= _GEN_34;
      end
    end else begin
      dst_d_r <= _GEN_34;
    end
    if (reset) begin // @[execute.scala 38:30]
      rcsr_id_r <= 12'h0; // @[execute.scala 38:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      rcsr_id_r <= io_rr2ex_rcsr_id; // @[execute.scala 97:21]
    end
    if (reset) begin // @[execute.scala 39:30]
      special_r <= 2'h0; // @[execute.scala 39:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      special_r <= io_rr2ex_special; // @[execute.scala 98:21]
    end
    if (reset) begin // @[execute.scala 40:30]
      alu64_r <= 1'h0; // @[execute.scala 40:30]
    end else if (hs_in) begin // @[execute.scala 70:26]
      alu64_r <= alu64;
    end
    if (reset) begin // @[execute.scala 41:30]
      indi_r <= 2'h0; // @[execute.scala 41:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      if (~memAlign) begin // @[execute.scala 105:24]
        indi_r <= 2'h0; // @[execute.scala 107:20]
      end else begin
        indi_r <= io_rr2ex_indi; // @[execute.scala 99:21]
      end
    end
    if (reset) begin // @[execute.scala 42:30]
      next_pc_r <= 64'h0; // @[execute.scala 42:30]
    end else if (hs_in) begin // @[execute.scala 170:16]
      if (_real_target_T) begin // @[Mux.scala 47:69]
        next_pc_r <= io_rr2ex_rs2_d;
      end else if (_real_target_T_1) begin // @[Mux.scala 47:69]
        next_pc_r <= _real_target_T_6;
      end else begin
        next_pc_r <= _real_target_T_10;
      end
    end else if (io_updateNextPc_valid) begin // @[execute.scala 78:32]
      next_pc_r <= io_updateNextPc_seq_pc; // @[execute.scala 79:19]
    end
    if (reset) begin // @[execute.scala 43:30]
      recov_r <= 1'h0; // @[execute.scala 43:30]
    end else if (hs_in) begin // @[execute.scala 86:16]
      recov_r <= _GEN_15;
    end
    if (reset) begin // @[execute.scala 44:30]
      valid_r <= 1'h0; // @[execute.scala 44:30]
    end else begin
      valid_r <= _GEN_59;
    end
    if (reset) begin // @[execute.scala 118:24]
      state <= 1'h0; // @[execute.scala 118:24]
    end else if (_io_rr2ex_stall_T) begin // @[execute.scala 127:26]
      if (state) begin // @[execute.scala 138:33]
        if (alu_io_valid) begin // @[execute.scala 139:31]
          state <= 1'h0; // @[execute.scala 140:29]
        end else begin
          state <= _GEN_49;
        end
      end else begin
        state <= _GEN_49;
      end
    end
    if (reset) begin // @[execute.scala 119:27]
      drop_alu <= 1'h0; // @[execute.scala 119:27]
    end else if (_io_rr2ex_stall_T) begin // @[execute.scala 127:26]
      if (state) begin // @[execute.scala 138:33]
        if (alu_io_valid) begin // @[execute.scala 139:31]
          drop_alu <= 1'h0; // @[execute.scala 143:29]
        end
      end
    end else begin
      drop_alu <= _GEN_58;
    end
    if (reset) begin // @[execute.scala 154:27]
      forceJmp_seq_pc <= 64'h0; // @[execute.scala 154:27]
    end else if (_T_2) begin // @[execute.scala 173:19]
      if (hs_in & ~io_rr2ex_excep_en & real_is_target & io_rr2ex_jmp_type != 2'h0) begin // @[execute.scala 174:92]
        if (_real_target_T) begin // @[Mux.scala 47:69]
          forceJmp_seq_pc <= io_rr2ex_rs2_d;
        end else begin
          forceJmp_seq_pc <= _real_target_T_11;
        end
      end
    end
    if (reset) begin // @[execute.scala 154:27]
      forceJmp_valid <= 1'h0; // @[execute.scala 154:27]
    end else begin
      forceJmp_valid <= _GEN_68;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  drop_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  stall_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  inst_r = _RAND_2[31:0];
  _RAND_3 = {2{`RANDOM}};
  pc_r = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  excep_r_cause = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  excep_r_tval = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  excep_r_en = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  excep_r_pc = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  excep_r_etype = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  ctrl_r_dcMode = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  ctrl_r_writeRegEn = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ctrl_r_writeCSREn = _RAND_11[0:0];
  _RAND_12 = {2{`RANDOM}};
  mem_addr_r = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  mem_data_r = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  csr_id_r = _RAND_14[11:0];
  _RAND_15 = {2{`RANDOM}};
  csr_d_r = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  dst_r = _RAND_16[4:0];
  _RAND_17 = {2{`RANDOM}};
  dst_d_r = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  rcsr_id_r = _RAND_18[11:0];
  _RAND_19 = {1{`RANDOM}};
  special_r = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  alu64_r = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  indi_r = _RAND_21[1:0];
  _RAND_22 = {2{`RANDOM}};
  next_pc_r = _RAND_22[63:0];
  _RAND_23 = {1{`RANDOM}};
  recov_r = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_r = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  state = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  drop_alu = _RAND_26[0:0];
  _RAND_27 = {2{`RANDOM}};
  forceJmp_seq_pc = _RAND_27[63:0];
  _RAND_28 = {1{`RANDOM}};
  forceJmp_valid = _RAND_28[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_Memory(
  input         clock,
  input         reset,
  input  [31:0] io_ex2mem_inst,
  input  [63:0] io_ex2mem_pc,
  input  [63:0] io_ex2mem_excep_cause,
  input  [63:0] io_ex2mem_excep_tval,
  input         io_ex2mem_excep_en,
  input  [63:0] io_ex2mem_excep_pc,
  input  [1:0]  io_ex2mem_excep_etype,
  input  [4:0]  io_ex2mem_ctrl_dcMode,
  input         io_ex2mem_ctrl_writeRegEn,
  input         io_ex2mem_ctrl_writeCSREn,
  input  [63:0] io_ex2mem_mem_addr,
  input  [63:0] io_ex2mem_mem_data,
  input  [11:0] io_ex2mem_csr_id,
  input  [63:0] io_ex2mem_csr_d,
  input  [4:0]  io_ex2mem_dst,
  input  [63:0] io_ex2mem_dst_d,
  input  [11:0] io_ex2mem_rcsr_id,
  input  [1:0]  io_ex2mem_special,
  input  [1:0]  io_ex2mem_indi,
  output        io_ex2mem_drop,
  output        io_ex2mem_stall,
  input         io_ex2mem_recov,
  input         io_ex2mem_valid,
  output        io_ex2mem_ready,
  output [31:0] io_mem2rb_inst,
  output [63:0] io_mem2rb_pc,
  output [63:0] io_mem2rb_excep_cause,
  output [63:0] io_mem2rb_excep_tval,
  output        io_mem2rb_excep_en,
  output [63:0] io_mem2rb_excep_pc,
  output [1:0]  io_mem2rb_excep_etype,
  output [11:0] io_mem2rb_csr_id,
  output [63:0] io_mem2rb_csr_d,
  output        io_mem2rb_csr_en,
  output [4:0]  io_mem2rb_dst,
  output [63:0] io_mem2rb_dst_d,
  output        io_mem2rb_dst_en,
  output [11:0] io_mem2rb_rcsr_id,
  output [1:0]  io_mem2rb_special,
  output        io_mem2rb_is_mmio,
  input         io_mem2rb_drop,
  input         io_mem2rb_stall,
  output        io_mem2rb_recov,
  output        io_mem2rb_valid,
  input         io_mem2rb_ready,
  output [31:0] io_dataRW_addr,
  input  [63:0] io_dataRW_rdata,
  input         io_dataRW_rvalid,
  output [63:0] io_dataRW_wdata,
  output [4:0]  io_dataRW_dc_mode,
  output [4:0]  io_dataRW_amo,
  input         io_dataRW_ready,
  output [63:0] io_va2pa_vaddr,
  output        io_va2pa_vvalid,
  output [1:0]  io_va2pa_m_type,
  input  [31:0] io_va2pa_paddr,
  input         io_va2pa_pvalid,
  input  [63:0] io_va2pa_tlb_excep_cause,
  input  [63:0] io_va2pa_tlb_excep_tval,
  input         io_va2pa_tlb_excep_en,
  output [4:0]  io_d_mem1_id,
  output [63:0] io_d_mem1_data,
  output [1:0]  io_d_mem1_state,
  output [4:0]  io_d_mem2_id,
  output [63:0] io_d_mem2_data,
  output [1:0]  io_d_mem2_state,
  output [4:0]  io_d_mem3_id,
  output [63:0] io_d_mem3_data,
  output [1:0]  io_d_mem3_state
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
`endif // RANDOMIZE_REG_INIT
  reg  drop2_r; // @[memory.scala 95:26]
  reg  stall2_r; // @[memory.scala 98:27]
  wire  drop2_in = drop2_r | io_mem2rb_drop; // @[memory.scala 103:31]
  wire  _stall3_in_T = ~io_mem2rb_drop; // @[memory.scala 105:34]
  wire  _stall1_in_T = ~drop2_in; // @[memory.scala 107:34]
  reg [31:0] inst1_r; // @[memory.scala 111:30]
  reg [63:0] pc1_r; // @[memory.scala 112:30]
  reg [63:0] excep1_r_cause; // @[memory.scala 113:30]
  reg [63:0] excep1_r_tval; // @[memory.scala 113:30]
  reg  excep1_r_en; // @[memory.scala 113:30]
  reg [63:0] excep1_r_pc; // @[memory.scala 113:30]
  reg [1:0] excep1_r_etype; // @[memory.scala 113:30]
  reg [4:0] ctrl1_r_dcMode; // @[memory.scala 114:30]
  reg [63:0] mem_addr1_r; // @[memory.scala 115:30]
  reg [63:0] mem_data1_r; // @[memory.scala 116:30]
  reg [4:0] dst1_r; // @[memory.scala 117:30]
  reg [63:0] dst_d1_r; // @[memory.scala 118:30]
  reg  dst_en1_r; // @[memory.scala 119:30]
  reg [11:0] csr_id1_r; // @[memory.scala 120:30]
  reg [63:0] csr_d1_r; // @[memory.scala 121:30]
  reg  csr_en1_r; // @[memory.scala 122:30]
  reg [11:0] rcsr_id1_r; // @[memory.scala 123:30]
  reg [1:0] special1_r; // @[memory.scala 124:30]
  reg [1:0] indi1_r; // @[memory.scala 125:30]
  reg  recov1_r; // @[memory.scala 126:30]
  reg  valid1_r; // @[memory.scala 128:30]
  reg  is_tlb_r; // @[memory.scala 134:30]
  reg  drop_tlb; // @[memory.scala 135:30]
  wire  hs_in = io_ex2mem_ready & io_ex2mem_valid; // @[memory.scala 137:35]
  wire [4:0] _GEN_10 = hs_in ? io_ex2mem_ctrl_dcMode : ctrl1_r_dcMode; // @[memory.scala 142:16 memory.scala 146:21 memory.scala 114:30]
  wire  access_tlb = io_ex2mem_ctrl_dcMode != 5'h0; // @[memory.scala 160:45]
  reg  valid2_r; // @[memory.scala 214:30]
  reg  valid3_r; // @[memory.scala 343:30]
  reg [4:0] ctrl2_r_dcMode; // @[memory.scala 201:30]
  wire  is_dc_r = ctrl2_r_dcMode != 5'h0; // @[memory.scala 254:39]
  wire  _dc_valid3_T = ~is_dc_r; // @[memory.scala 367:21]
  reg  drop_dc; // @[memory.scala 255:30]
  wire  dc_valid3 = ~is_dc_r | io_dataRW_rvalid & ~drop_dc; // @[memory.scala 367:30]
  wire  _T_34 = valid2_r & dc_valid3; // @[memory.scala 370:29]
  wire  _GEN_167 = valid3_r & ~io_mem2rb_ready ? 1'h0 : _T_34; // @[memory.scala 369:34 memory.scala 141:25]
  wire  hs2 = _stall3_in_T & _GEN_167; // @[memory.scala 368:20 memory.scala 141:25]
  wire  inp_tlb_valid2 = io_va2pa_pvalid | io_va2pa_tlb_excep_en; // @[memory.scala 260:42]
  wire  _tlb_valid2_T_1 = ~drop_tlb; // @[memory.scala 282:55]
  wire  tlb_valid2 = ~is_tlb_r | inp_tlb_valid2 & ~drop_tlb; // @[memory.scala 282:33]
  wire  _T_23 = valid1_r & tlb_valid2; // @[memory.scala 289:29]
  wire  _GEN_89 = valid2_r & ~hs2 ? 1'h0 : _T_23; // @[memory.scala 288:31 memory.scala 141:9]
  wire  hs1 = _stall1_in_T & _GEN_89; // @[memory.scala 287:20 memory.scala 141:9]
  wire  _io_va2pa_vvalid_T_2 = ~hs1; // @[memory.scala 162:49]
  wire  _GEN_26 = valid1_r & _io_va2pa_vvalid_T_2 ? 1'h0 : io_ex2mem_valid; // @[memory.scala 167:31 memory.scala 165:21]
  wire  _GEN_28 = hs1 ? 1'h0 : valid1_r; // @[memory.scala 177:24 memory.scala 178:22 memory.scala 128:30]
  wire  _GEN_29 = hs1 ? 1'h0 : is_tlb_r; // @[memory.scala 177:24 memory.scala 179:22 memory.scala 134:30]
  wire  _GEN_30 = hs_in | _GEN_28; // @[memory.scala 173:20 memory.scala 174:22]
  wire  _GEN_31 = hs_in ? access_tlb : _GEN_29; // @[memory.scala 173:20 memory.scala 175:22]
  wire  _GEN_32 = hs_in ? access_tlb : _stall1_in_T & is_tlb_r & ~hs1; // @[memory.scala 173:20 memory.scala 176:29 memory.scala 162:21]
  wire  _GEN_33 = _stall1_in_T & _GEN_30; // @[memory.scala 172:20 memory.scala 182:18]
  wire  _GEN_34 = _stall1_in_T & _GEN_31; // @[memory.scala 172:20 memory.scala 184:18]
  wire [1:0] _GEN_37 = valid1_r ? 2'h2 : 2'h0; // @[memory.scala 192:25 memory.scala 193:25 memory.scala 195:25]
  wire [1:0] _GEN_38 = valid1_r & ~(ctrl1_r_dcMode[2] | indi1_r[1]) ? 2'h1 : _GEN_37; // @[memory.scala 190:80 memory.scala 191:25]
  reg [31:0] inst2_r; // @[memory.scala 198:30]
  reg [63:0] pc2_r; // @[memory.scala 199:30]
  reg [63:0] excep2_r_cause; // @[memory.scala 200:30]
  reg [63:0] excep2_r_tval; // @[memory.scala 200:30]
  reg  excep2_r_en; // @[memory.scala 200:30]
  reg [63:0] excep2_r_pc; // @[memory.scala 200:30]
  reg [1:0] excep2_r_etype; // @[memory.scala 200:30]
  reg [63:0] mem_data2_r; // @[memory.scala 202:30]
  reg [4:0] dst2_r; // @[memory.scala 203:30]
  reg [63:0] dst_d2_r; // @[memory.scala 204:30]
  reg  dst_en2_r; // @[memory.scala 205:30]
  reg [11:0] csr_id2_r; // @[memory.scala 206:30]
  reg [63:0] csr_d2_r; // @[memory.scala 207:30]
  reg  csr_en2_r; // @[memory.scala 208:30]
  reg [11:0] rcsr_id2_r; // @[memory.scala 209:30]
  reg [1:0] special2_r; // @[memory.scala 210:30]
  reg [31:0] paddr2_r; // @[memory.scala 211:30]
  reg  recov2_r; // @[memory.scala 213:30]
  reg  dc_hs_r; // @[memory.scala 215:30]
  reg [31:0] lr_addr_r; // @[memory.scala 217:30]
  reg  lr_valid_r; // @[memory.scala 218:30]
  wire  stage2_is_excep = excep1_r_en | io_va2pa_tlb_excep_en; // @[memory.scala 227:39]
  wire  _GEN_41 = indi1_r[0] & ~stage2_is_excep | lr_valid_r; // @[memory.scala 245:55 memory.scala 246:25 memory.scala 218:30]
  wire [1:0] _GEN_46 = hs1 ? excep1_r_etype : excep2_r_etype; // @[memory.scala 228:14 memory.scala 231:21 memory.scala 200:30]
  wire [63:0] _GEN_47 = hs1 ? excep1_r_pc : excep2_r_pc; // @[memory.scala 228:14 memory.scala 231:21 memory.scala 200:30]
  wire  _GEN_48 = hs1 ? excep1_r_en : excep2_r_en; // @[memory.scala 228:14 memory.scala 231:21 memory.scala 200:30]
  wire [63:0] _GEN_49 = hs1 ? excep1_r_tval : excep2_r_tval; // @[memory.scala 228:14 memory.scala 231:21 memory.scala 200:30]
  wire [63:0] _GEN_50 = hs1 ? excep1_r_cause : excep2_r_cause; // @[memory.scala 228:14 memory.scala 231:21 memory.scala 200:30]
  wire [4:0] _GEN_55 = hs1 ? ctrl1_r_dcMode : ctrl2_r_dcMode; // @[memory.scala 228:14 memory.scala 233:21 memory.scala 201:30]
  wire [63:0] _GEN_59 = hs1 ? dst_d1_r : dst_d2_r; // @[memory.scala 228:14 memory.scala 235:21 memory.scala 204:30]
  wire  _GEN_60 = hs1 ? dst_en1_r : dst_en2_r; // @[memory.scala 228:14 memory.scala 236:21 memory.scala 205:30]
  wire  _GEN_63 = hs1 ? csr_en1_r : csr_en2_r; // @[memory.scala 228:14 memory.scala 239:21 memory.scala 208:30]
  wire  _GEN_67 = hs1 ? recov1_r : recov2_r; // @[memory.scala 228:14 memory.scala 243:21 memory.scala 213:30]
  wire  sc_valid = io_va2pa_paddr == lr_addr_r & lr_valid_r; // @[memory.scala 261:52]
  wire [4:0] _GEN_71 = indi1_r[1] ? 5'h0 : ctrl1_r_dcMode; // @[memory.scala 270:41 memory.scala 271:31 memory.scala 276:31]
  wire [4:0] _GEN_72 = indi1_r[1] ? 5'h0 : _GEN_55; // @[memory.scala 270:41 memory.scala 272:29]
  wire  _GEN_73 = indi1_r[1] | _GEN_60; // @[memory.scala 270:41 memory.scala 273:25]
  wire [63:0] _GEN_74 = indi1_r[1] ? 64'h1 : _GEN_59; // @[memory.scala 270:41 memory.scala 274:25]
  wire [4:0] _GEN_75 = indi1_r[1] & sc_valid ? ctrl1_r_dcMode : _GEN_71; // @[memory.scala 266:53 memory.scala 267:31]
  wire  _GEN_76 = indi1_r[1] & sc_valid | _GEN_73; // @[memory.scala 266:53 memory.scala 268:25]
  wire [4:0] _GEN_78 = indi1_r[1] & sc_valid ? _GEN_55 : _GEN_72; // @[memory.scala 266:53]
  wire [4:0] _GEN_79 = stage2_is_excep ? 5'h0 : _GEN_75; // @[memory.scala 263:30 memory.scala 264:31]
  wire [4:0] _GEN_80 = stage2_is_excep ? 5'h0 : _GEN_78; // @[memory.scala 263:30 memory.scala 265:29]
  wire  _GEN_81 = stage2_is_excep ? _GEN_60 : _GEN_76; // @[memory.scala 263:30]
  wire [4:0] _io_dataRW_dc_mode_T_2 = valid2_r & ~dc_hs_r ? ctrl2_r_dcMode : 5'h0; // @[memory.scala 279:33]
  wire [4:0] _GEN_84 = hs1 ? _GEN_80 : _GEN_55; // @[memory.scala 262:14]
  wire  _GEN_85 = hs1 ? _GEN_81 : _GEN_60; // @[memory.scala 262:14]
  wire  dc_hs = io_dataRW_dc_mode != 5'h0 & io_dataRW_ready; // @[memory.scala 283:48]
  wire  _GEN_87 = dc_hs | dc_hs_r; // @[memory.scala 284:16 memory.scala 285:17 memory.scala 215:30]
  wire  _T_26 = io_va2pa_tlb_excep_en & _tlb_valid2_T_1; // @[memory.scala 296:40]
  wire  _GEN_91 = ctrl1_r_dcMode != 5'h0 ? dc_hs : _GEN_87; // @[memory.scala 306:52 memory.scala 307:25]
  wire  _GEN_94 = io_va2pa_tlb_excep_en & _tlb_valid2_T_1 | _GEN_48; // @[memory.scala 296:53 memory.scala 299:33]
  wire  _GEN_106 = io_va2pa_tlb_excep_en & _tlb_valid2_T_1 | _GEN_67; // @[memory.scala 296:53 memory.scala 221:57]
  wire  _GEN_108 = hs2 ? 1'h0 : valid2_r; // @[memory.scala 309:24 memory.scala 310:22 memory.scala 214:30]
  wire  _GEN_110 = hs1 | _GEN_108; // @[memory.scala 294:18 memory.scala 295:22]
  wire  _GEN_124 = hs1 & _T_26; // @[memory.scala 294:18 memory.scala 100:13]
  wire  _GEN_127 = _stall3_in_T & _GEN_110; // @[memory.scala 293:20 memory.scala 314:18]
  wire  _GEN_141 = _stall3_in_T & _GEN_124; // @[memory.scala 293:20 memory.scala 100:13]
  wire [1:0] _GEN_145 = valid2_r ? 2'h2 : 2'h0; // @[memory.scala 324:25 memory.scala 325:25 memory.scala 327:25]
  wire [1:0] _GEN_146 = valid2_r & _dc_valid3_T ? 2'h1 : _GEN_145; // @[memory.scala 322:37 memory.scala 323:25]
  reg [31:0] inst3_r; // @[memory.scala 330:30]
  reg [63:0] pc3_r; // @[memory.scala 331:30]
  reg [63:0] excep3_r_cause; // @[memory.scala 332:30]
  reg [63:0] excep3_r_tval; // @[memory.scala 332:30]
  reg  excep3_r_en; // @[memory.scala 332:30]
  reg [63:0] excep3_r_pc; // @[memory.scala 332:30]
  reg [1:0] excep3_r_etype; // @[memory.scala 332:30]
  reg [4:0] dst3_r; // @[memory.scala 333:30]
  reg [63:0] dst_d3_r; // @[memory.scala 334:30]
  reg  dst_en3_r; // @[memory.scala 335:30]
  reg [11:0] csr_id3_r; // @[memory.scala 336:30]
  reg [63:0] csr_d3_r; // @[memory.scala 337:30]
  reg  csr_en3_r; // @[memory.scala 338:30]
  reg [11:0] rcsr_id3_r; // @[memory.scala 339:30]
  reg [1:0] special3_r; // @[memory.scala 340:30]
  reg  is_mmio_r; // @[memory.scala 341:30]
  reg  recov3_r; // @[memory.scala 342:30]
  wire [63:0] _GEN_156 = hs2 ? dst_d2_r : dst_d3_r; // @[memory.scala 349:14 memory.scala 354:21 memory.scala 334:30]
  wire  _GEN_170 = io_mem2rb_ready ? 1'h0 : valid3_r; // @[memory.scala 380:27 memory.scala 381:22 memory.scala 343:30]
  wire  _GEN_171 = hs2 | _GEN_170; // @[memory.scala 375:19 memory.scala 376:22]
  wire  _GEN_173 = _stall3_in_T & _GEN_171; // @[memory.scala 374:26 memory.scala 384:18]
  assign io_ex2mem_drop = drop2_r | io_mem2rb_drop; // @[memory.scala 103:31]
  assign io_ex2mem_stall = stall2_r & _stall3_in_T | io_mem2rb_stall; // @[memory.scala 106:45]
  assign io_ex2mem_ready = _stall1_in_T & _GEN_26; // @[memory.scala 166:20 memory.scala 165:21]
  assign io_mem2rb_inst = inst3_r; // @[memory.scala 386:25]
  assign io_mem2rb_pc = pc3_r; // @[memory.scala 387:25]
  assign io_mem2rb_excep_cause = excep3_r_cause; // @[memory.scala 388:25]
  assign io_mem2rb_excep_tval = excep3_r_tval; // @[memory.scala 388:25]
  assign io_mem2rb_excep_en = excep3_r_en; // @[memory.scala 388:25]
  assign io_mem2rb_excep_pc = excep3_r_pc; // @[memory.scala 388:25]
  assign io_mem2rb_excep_etype = excep3_r_etype; // @[memory.scala 388:25]
  assign io_mem2rb_csr_id = csr_id3_r; // @[memory.scala 389:25]
  assign io_mem2rb_csr_d = csr_d3_r; // @[memory.scala 390:25]
  assign io_mem2rb_csr_en = csr_en3_r; // @[memory.scala 391:25]
  assign io_mem2rb_dst = dst3_r; // @[memory.scala 392:25]
  assign io_mem2rb_dst_d = dst_d3_r; // @[memory.scala 393:25]
  assign io_mem2rb_dst_en = dst_en3_r; // @[memory.scala 394:25]
  assign io_mem2rb_rcsr_id = rcsr_id3_r; // @[memory.scala 395:25]
  assign io_mem2rb_special = special3_r; // @[memory.scala 396:25]
  assign io_mem2rb_is_mmio = is_mmio_r; // @[memory.scala 397:25]
  assign io_mem2rb_recov = recov3_r; // @[memory.scala 398:25]
  assign io_mem2rb_valid = valid3_r; // @[memory.scala 399:25]
  assign io_dataRW_addr = hs1 ? io_va2pa_paddr : paddr2_r; // @[memory.scala 257:29]
  assign io_dataRW_wdata = hs1 ? mem_data1_r : mem_data2_r; // @[memory.scala 258:29]
  assign io_dataRW_dc_mode = hs1 ? _GEN_79 : _io_dataRW_dc_mode_T_2; // @[memory.scala 262:14 memory.scala 279:27]
  assign io_dataRW_amo = hs1 ? inst1_r[31:27] : inst2_r[31:27]; // @[memory.scala 259:29]
  assign io_va2pa_vaddr = hs_in ? io_ex2mem_mem_addr : mem_addr1_r; // @[memory.scala 161:27]
  assign io_va2pa_vvalid = _stall1_in_T ? _GEN_32 : _stall1_in_T & is_tlb_r & ~hs1; // @[memory.scala 172:20 memory.scala 162:21]
  assign io_va2pa_m_type = _GEN_10[3] ? 2'h3 : 2'h2; // @[memory.scala 164:27]
  assign io_d_mem1_id = dst1_r; // @[memory.scala 186:20]
  assign io_d_mem1_data = dst_d1_r; // @[memory.scala 187:20]
  assign io_d_mem1_state = ~dst_en1_r ? 2'h0 : _GEN_38; // @[memory.scala 188:21 memory.scala 189:25]
  assign io_d_mem2_id = dst2_r; // @[memory.scala 318:20]
  assign io_d_mem2_data = dst_d2_r; // @[memory.scala 319:20]
  assign io_d_mem2_state = ~dst_en2_r ? 2'h0 : _GEN_146; // @[memory.scala 320:21 memory.scala 321:25]
  assign io_d_mem3_id = dst3_r; // @[memory.scala 401:20]
  assign io_d_mem3_data = dst_d3_r; // @[memory.scala 402:20]
  assign io_d_mem3_state = valid3_r & dst_en3_r ? 2'h1 : 2'h0; // @[memory.scala 403:32 memory.scala 404:25 memory.scala 406:25]
  always @(posedge clock) begin
    if (reset) begin // @[memory.scala 95:26]
      drop2_r <= 1'h0; // @[memory.scala 95:26]
    end else begin
      drop2_r <= _GEN_141;
    end
    if (reset) begin // @[memory.scala 98:27]
      stall2_r <= 1'h0; // @[memory.scala 98:27]
    end else begin
      stall2_r <= _GEN_141;
    end
    if (reset) begin // @[memory.scala 111:30]
      inst1_r <= 32'h0; // @[memory.scala 111:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      inst1_r <= io_ex2mem_inst; // @[memory.scala 143:21]
    end
    if (reset) begin // @[memory.scala 112:30]
      pc1_r <= 64'h0; // @[memory.scala 112:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      pc1_r <= io_ex2mem_pc; // @[memory.scala 144:21]
    end
    if (reset) begin // @[memory.scala 113:30]
      excep1_r_cause <= 64'h0; // @[memory.scala 113:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      excep1_r_cause <= io_ex2mem_excep_cause; // @[memory.scala 145:21]
    end
    if (reset) begin // @[memory.scala 113:30]
      excep1_r_tval <= 64'h0; // @[memory.scala 113:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      excep1_r_tval <= io_ex2mem_excep_tval; // @[memory.scala 145:21]
    end
    if (reset) begin // @[memory.scala 113:30]
      excep1_r_en <= 1'h0; // @[memory.scala 113:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      excep1_r_en <= io_ex2mem_excep_en; // @[memory.scala 145:21]
    end
    if (reset) begin // @[memory.scala 113:30]
      excep1_r_pc <= 64'h0; // @[memory.scala 113:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      excep1_r_pc <= io_ex2mem_excep_pc; // @[memory.scala 145:21]
    end
    if (reset) begin // @[memory.scala 113:30]
      excep1_r_etype <= 2'h0; // @[memory.scala 113:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      excep1_r_etype <= io_ex2mem_excep_etype; // @[memory.scala 145:21]
    end
    if (reset) begin // @[memory.scala 114:30]
      ctrl1_r_dcMode <= 5'h0; // @[memory.scala 114:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      ctrl1_r_dcMode <= io_ex2mem_ctrl_dcMode; // @[memory.scala 146:21]
    end
    if (reset) begin // @[memory.scala 115:30]
      mem_addr1_r <= 64'h0; // @[memory.scala 115:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      mem_addr1_r <= io_ex2mem_mem_addr; // @[memory.scala 147:21]
    end
    if (reset) begin // @[memory.scala 116:30]
      mem_data1_r <= 64'h0; // @[memory.scala 116:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      mem_data1_r <= io_ex2mem_mem_data; // @[memory.scala 148:21]
    end
    if (reset) begin // @[memory.scala 117:30]
      dst1_r <= 5'h0; // @[memory.scala 117:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      dst1_r <= io_ex2mem_dst; // @[memory.scala 149:21]
    end
    if (reset) begin // @[memory.scala 118:30]
      dst_d1_r <= 64'h0; // @[memory.scala 118:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      dst_d1_r <= io_ex2mem_dst_d; // @[memory.scala 150:21]
    end
    if (reset) begin // @[memory.scala 119:30]
      dst_en1_r <= 1'h0; // @[memory.scala 119:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      dst_en1_r <= io_ex2mem_ctrl_writeRegEn; // @[memory.scala 151:21]
    end
    if (reset) begin // @[memory.scala 120:30]
      csr_id1_r <= 12'h0; // @[memory.scala 120:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      csr_id1_r <= io_ex2mem_csr_id; // @[memory.scala 152:21]
    end
    if (reset) begin // @[memory.scala 121:30]
      csr_d1_r <= 64'h0; // @[memory.scala 121:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      csr_d1_r <= io_ex2mem_csr_d; // @[memory.scala 153:21]
    end
    if (reset) begin // @[memory.scala 122:30]
      csr_en1_r <= 1'h0; // @[memory.scala 122:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      csr_en1_r <= io_ex2mem_ctrl_writeCSREn; // @[memory.scala 154:21]
    end
    if (reset) begin // @[memory.scala 123:30]
      rcsr_id1_r <= 12'h0; // @[memory.scala 123:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      rcsr_id1_r <= io_ex2mem_rcsr_id; // @[memory.scala 155:21]
    end
    if (reset) begin // @[memory.scala 124:30]
      special1_r <= 2'h0; // @[memory.scala 124:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      special1_r <= io_ex2mem_special; // @[memory.scala 157:21]
    end
    if (reset) begin // @[memory.scala 125:30]
      indi1_r <= 2'h0; // @[memory.scala 125:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      indi1_r <= io_ex2mem_indi; // @[memory.scala 156:21]
    end
    if (reset) begin // @[memory.scala 126:30]
      recov1_r <= 1'h0; // @[memory.scala 126:30]
    end else if (hs_in) begin // @[memory.scala 142:16]
      recov1_r <= io_ex2mem_recov; // @[memory.scala 158:21]
    end
    if (reset) begin // @[memory.scala 128:30]
      valid1_r <= 1'h0; // @[memory.scala 128:30]
    end else begin
      valid1_r <= _GEN_33;
    end
    if (reset) begin // @[memory.scala 134:30]
      is_tlb_r <= 1'h0; // @[memory.scala 134:30]
    end else begin
      is_tlb_r <= _GEN_34;
    end
    if (reset) begin // @[memory.scala 135:30]
      drop_tlb <= 1'h0; // @[memory.scala 135:30]
    end else if (inp_tlb_valid2 & drop_tlb) begin // @[memory.scala 224:65]
      drop_tlb <= 1'h0; // @[memory.scala 225:18]
    end else if (!(_stall1_in_T)) begin // @[memory.scala 172:20]
      drop_tlb <= is_tlb_r & ~io_va2pa_pvalid; // @[memory.scala 183:18]
    end
    if (reset) begin // @[memory.scala 214:30]
      valid2_r <= 1'h0; // @[memory.scala 214:30]
    end else begin
      valid2_r <= _GEN_127;
    end
    if (reset) begin // @[memory.scala 343:30]
      valid3_r <= 1'h0; // @[memory.scala 343:30]
    end else begin
      valid3_r <= _GEN_173;
    end
    if (reset) begin // @[memory.scala 201:30]
      ctrl2_r_dcMode <= 5'h0; // @[memory.scala 201:30]
    end else if (_stall3_in_T) begin // @[memory.scala 293:20]
      if (hs1) begin // @[memory.scala 294:18]
        if (io_va2pa_tlb_excep_en & _tlb_valid2_T_1) begin // @[memory.scala 296:53]
          ctrl2_r_dcMode <= 5'h0; // @[memory.scala 302:29]
        end else begin
          ctrl2_r_dcMode <= _GEN_84;
        end
      end else begin
        ctrl2_r_dcMode <= _GEN_84;
      end
    end else begin
      ctrl2_r_dcMode <= _GEN_84;
    end
    if (reset) begin // @[memory.scala 255:30]
      drop_dc <= 1'h0; // @[memory.scala 255:30]
    end else if (io_dataRW_rvalid) begin // @[memory.scala 364:27]
      drop_dc <= 1'h0; // @[memory.scala 365:17]
    end else if (!(_stall3_in_T)) begin // @[memory.scala 293:20]
      drop_dc <= is_dc_r & ~io_dataRW_rvalid; // @[memory.scala 315:18]
    end
    if (reset) begin // @[memory.scala 198:30]
      inst2_r <= 32'h0; // @[memory.scala 198:30]
    end else if (hs1) begin // @[memory.scala 228:14]
      inst2_r <= inst1_r; // @[memory.scala 229:21]
    end
    if (reset) begin // @[memory.scala 199:30]
      pc2_r <= 64'h0; // @[memory.scala 199:30]
    end else if (hs1) begin // @[memory.scala 228:14]
      pc2_r <= pc1_r; // @[memory.scala 230:21]
    end
    if (reset) begin // @[memory.scala 200:30]
      excep2_r_cause <= 64'h0; // @[memory.scala 200:30]
    end else if (_stall3_in_T) begin // @[memory.scala 293:20]
      if (hs1) begin // @[memory.scala 294:18]
        if (io_va2pa_tlb_excep_en & _tlb_valid2_T_1) begin // @[memory.scala 296:53]
          excep2_r_cause <= io_va2pa_tlb_excep_cause; // @[memory.scala 297:33]
        end else begin
          excep2_r_cause <= _GEN_50;
        end
      end else begin
        excep2_r_cause <= _GEN_50;
      end
    end else begin
      excep2_r_cause <= _GEN_50;
    end
    if (reset) begin // @[memory.scala 200:30]
      excep2_r_tval <= 64'h0; // @[memory.scala 200:30]
    end else if (_stall3_in_T) begin // @[memory.scala 293:20]
      if (hs1) begin // @[memory.scala 294:18]
        if (io_va2pa_tlb_excep_en & _tlb_valid2_T_1) begin // @[memory.scala 296:53]
          excep2_r_tval <= io_va2pa_tlb_excep_tval; // @[memory.scala 298:33]
        end else begin
          excep2_r_tval <= _GEN_49;
        end
      end else begin
        excep2_r_tval <= _GEN_49;
      end
    end else begin
      excep2_r_tval <= _GEN_49;
    end
    if (reset) begin // @[memory.scala 200:30]
      excep2_r_en <= 1'h0; // @[memory.scala 200:30]
    end else if (_stall3_in_T) begin // @[memory.scala 293:20]
      if (hs1) begin // @[memory.scala 294:18]
        excep2_r_en <= _GEN_94;
      end else begin
        excep2_r_en <= _GEN_48;
      end
    end else begin
      excep2_r_en <= _GEN_48;
    end
    if (reset) begin // @[memory.scala 200:30]
      excep2_r_pc <= 64'h0; // @[memory.scala 200:30]
    end else if (_stall3_in_T) begin // @[memory.scala 293:20]
      if (hs1) begin // @[memory.scala 294:18]
        if (io_va2pa_tlb_excep_en & _tlb_valid2_T_1) begin // @[memory.scala 296:53]
          excep2_r_pc <= pc1_r; // @[memory.scala 300:33]
        end else begin
          excep2_r_pc <= _GEN_47;
        end
      end else begin
        excep2_r_pc <= _GEN_47;
      end
    end else begin
      excep2_r_pc <= _GEN_47;
    end
    if (reset) begin // @[memory.scala 200:30]
      excep2_r_etype <= 2'h0; // @[memory.scala 200:30]
    end else if (_stall3_in_T) begin // @[memory.scala 293:20]
      if (hs1) begin // @[memory.scala 294:18]
        if (io_va2pa_tlb_excep_en & _tlb_valid2_T_1) begin // @[memory.scala 296:53]
          excep2_r_etype <= 2'h0; // @[memory.scala 301:33]
        end else begin
          excep2_r_etype <= _GEN_46;
        end
      end else begin
        excep2_r_etype <= _GEN_46;
      end
    end else begin
      excep2_r_etype <= _GEN_46;
    end
    if (reset) begin // @[memory.scala 202:30]
      mem_data2_r <= 64'h0; // @[memory.scala 202:30]
    end else if (hs1) begin // @[memory.scala 228:14]
      mem_data2_r <= mem_data1_r; // @[memory.scala 232:21]
    end
    if (reset) begin // @[memory.scala 203:30]
      dst2_r <= 5'h0; // @[memory.scala 203:30]
    end else if (hs1) begin // @[memory.scala 228:14]
      dst2_r <= dst1_r; // @[memory.scala 234:21]
    end
    if (reset) begin // @[memory.scala 204:30]
      dst_d2_r <= 64'h0; // @[memory.scala 204:30]
    end else if (hs1) begin // @[memory.scala 262:14]
      if (stage2_is_excep) begin // @[memory.scala 263:30]
        dst_d2_r <= _GEN_59;
      end else if (indi1_r[1] & sc_valid) begin // @[memory.scala 266:53]
        dst_d2_r <= 64'h0; // @[memory.scala 269:25]
      end else begin
        dst_d2_r <= _GEN_74;
      end
    end else begin
      dst_d2_r <= _GEN_59;
    end
    if (reset) begin // @[memory.scala 205:30]
      dst_en2_r <= 1'h0; // @[memory.scala 205:30]
    end else if (_stall3_in_T) begin // @[memory.scala 293:20]
      if (hs1) begin // @[memory.scala 294:18]
        if (io_va2pa_tlb_excep_en & _tlb_valid2_T_1) begin // @[memory.scala 296:53]
          dst_en2_r <= 1'h0; // @[memory.scala 303:29]
        end else begin
          dst_en2_r <= _GEN_85;
        end
      end else begin
        dst_en2_r <= _GEN_85;
      end
    end else begin
      dst_en2_r <= _GEN_85;
    end
    if (reset) begin // @[memory.scala 206:30]
      csr_id2_r <= 12'h0; // @[memory.scala 206:30]
    end else if (hs1) begin // @[memory.scala 228:14]
      csr_id2_r <= csr_id1_r; // @[memory.scala 237:21]
    end
    if (reset) begin // @[memory.scala 207:30]
      csr_d2_r <= 64'h0; // @[memory.scala 207:30]
    end else if (hs1) begin // @[memory.scala 228:14]
      csr_d2_r <= csr_d1_r; // @[memory.scala 238:21]
    end
    if (reset) begin // @[memory.scala 208:30]
      csr_en2_r <= 1'h0; // @[memory.scala 208:30]
    end else if (_stall3_in_T) begin // @[memory.scala 293:20]
      if (hs1) begin // @[memory.scala 294:18]
        if (io_va2pa_tlb_excep_en & _tlb_valid2_T_1) begin // @[memory.scala 296:53]
          csr_en2_r <= 1'h0; // @[memory.scala 304:29]
        end else begin
          csr_en2_r <= _GEN_63;
        end
      end else begin
        csr_en2_r <= _GEN_63;
      end
    end else begin
      csr_en2_r <= _GEN_63;
    end
    if (reset) begin // @[memory.scala 209:30]
      rcsr_id2_r <= 12'h0; // @[memory.scala 209:30]
    end else if (hs1) begin // @[memory.scala 228:14]
      rcsr_id2_r <= rcsr_id1_r; // @[memory.scala 240:21]
    end
    if (reset) begin // @[memory.scala 210:30]
      special2_r <= 2'h0; // @[memory.scala 210:30]
    end else if (hs1) begin // @[memory.scala 228:14]
      special2_r <= special1_r; // @[memory.scala 241:21]
    end
    if (reset) begin // @[memory.scala 211:30]
      paddr2_r <= 32'h0; // @[memory.scala 211:30]
    end else if (hs1) begin // @[memory.scala 228:14]
      paddr2_r <= io_va2pa_paddr; // @[memory.scala 244:21]
    end
    if (reset) begin // @[memory.scala 213:30]
      recov2_r <= 1'h0; // @[memory.scala 213:30]
    end else if (_stall3_in_T) begin // @[memory.scala 293:20]
      if (hs1) begin // @[memory.scala 294:18]
        recov2_r <= _GEN_106;
      end else begin
        recov2_r <= _GEN_67;
      end
    end else begin
      recov2_r <= _GEN_67;
    end
    if (reset) begin // @[memory.scala 215:30]
      dc_hs_r <= 1'h0; // @[memory.scala 215:30]
    end else if (_stall3_in_T) begin // @[memory.scala 293:20]
      if (hs1) begin // @[memory.scala 294:18]
        if (io_va2pa_tlb_excep_en & _tlb_valid2_T_1) begin // @[memory.scala 296:53]
          dc_hs_r <= _GEN_87;
        end else begin
          dc_hs_r <= _GEN_91;
        end
      end else if (hs2) begin // @[memory.scala 309:24]
        dc_hs_r <= 1'h0; // @[memory.scala 311:22]
      end else begin
        dc_hs_r <= _GEN_87;
      end
    end else begin
      dc_hs_r <= _GEN_87;
    end
    if (reset) begin // @[memory.scala 217:30]
      lr_addr_r <= 32'h0; // @[memory.scala 217:30]
    end else if (hs1) begin // @[memory.scala 228:14]
      if (indi1_r[0] & ~stage2_is_excep) begin // @[memory.scala 245:55]
        lr_addr_r <= io_va2pa_paddr; // @[memory.scala 247:25]
      end
    end
    if (reset) begin // @[memory.scala 218:30]
      lr_valid_r <= 1'h0; // @[memory.scala 218:30]
    end else if (hs1) begin // @[memory.scala 228:14]
      if (excep1_r_en & excep1_r_cause[63]) begin // @[memory.scala 249:48]
        lr_valid_r <= 1'h0; // @[memory.scala 250:25]
      end else begin
        lr_valid_r <= _GEN_41;
      end
    end
    if (reset) begin // @[memory.scala 330:30]
      inst3_r <= 32'h0; // @[memory.scala 330:30]
    end else if (hs2) begin // @[memory.scala 349:14]
      inst3_r <= inst2_r; // @[memory.scala 350:21]
    end
    if (reset) begin // @[memory.scala 331:30]
      pc3_r <= 64'h0; // @[memory.scala 331:30]
    end else if (hs2) begin // @[memory.scala 349:14]
      pc3_r <= pc2_r; // @[memory.scala 351:21]
    end
    if (reset) begin // @[memory.scala 332:30]
      excep3_r_cause <= 64'h0; // @[memory.scala 332:30]
    end else if (hs2) begin // @[memory.scala 349:14]
      excep3_r_cause <= excep2_r_cause; // @[memory.scala 352:21]
    end
    if (reset) begin // @[memory.scala 332:30]
      excep3_r_tval <= 64'h0; // @[memory.scala 332:30]
    end else if (hs2) begin // @[memory.scala 349:14]
      excep3_r_tval <= excep2_r_tval; // @[memory.scala 352:21]
    end
    if (reset) begin // @[memory.scala 332:30]
      excep3_r_en <= 1'h0; // @[memory.scala 332:30]
    end else if (hs2) begin // @[memory.scala 349:14]
      excep3_r_en <= excep2_r_en; // @[memory.scala 352:21]
    end
    if (reset) begin // @[memory.scala 332:30]
      excep3_r_pc <= 64'h0; // @[memory.scala 332:30]
    end else if (hs2) begin // @[memory.scala 349:14]
      excep3_r_pc <= excep2_r_pc; // @[memory.scala 352:21]
    end
    if (reset) begin // @[memory.scala 332:30]
      excep3_r_etype <= 2'h0; // @[memory.scala 332:30]
    end else if (hs2) begin // @[memory.scala 349:14]
      excep3_r_etype <= excep2_r_etype; // @[memory.scala 352:21]
    end
    if (reset) begin // @[memory.scala 333:30]
      dst3_r <= 5'h0; // @[memory.scala 333:30]
    end else if (hs2) begin // @[memory.scala 349:14]
      dst3_r <= dst2_r; // @[memory.scala 353:21]
    end
    if (reset) begin // @[memory.scala 334:30]
      dst_d3_r <= 64'h0; // @[memory.scala 334:30]
    end else if (_stall3_in_T) begin // @[memory.scala 374:26]
      if (hs2) begin // @[memory.scala 375:19]
        if (is_dc_r) begin // @[memory.scala 377:26]
          dst_d3_r <= io_dataRW_rdata; // @[memory.scala 378:26]
        end else begin
          dst_d3_r <= _GEN_156;
        end
      end else begin
        dst_d3_r <= _GEN_156;
      end
    end else begin
      dst_d3_r <= _GEN_156;
    end
    if (reset) begin // @[memory.scala 335:30]
      dst_en3_r <= 1'h0; // @[memory.scala 335:30]
    end else if (hs2) begin // @[memory.scala 349:14]
      dst_en3_r <= dst_en2_r; // @[memory.scala 355:21]
    end
    if (reset) begin // @[memory.scala 336:30]
      csr_id3_r <= 12'h0; // @[memory.scala 336:30]
    end else if (hs2) begin // @[memory.scala 349:14]
      csr_id3_r <= csr_id2_r; // @[memory.scala 356:21]
    end
    if (reset) begin // @[memory.scala 337:30]
      csr_d3_r <= 64'h0; // @[memory.scala 337:30]
    end else if (hs2) begin // @[memory.scala 349:14]
      csr_d3_r <= csr_d2_r; // @[memory.scala 357:21]
    end
    if (reset) begin // @[memory.scala 338:30]
      csr_en3_r <= 1'h0; // @[memory.scala 338:30]
    end else if (hs2) begin // @[memory.scala 349:14]
      csr_en3_r <= csr_en2_r; // @[memory.scala 358:21]
    end
    if (reset) begin // @[memory.scala 339:30]
      rcsr_id3_r <= 12'h0; // @[memory.scala 339:30]
    end else if (hs2) begin // @[memory.scala 349:14]
      rcsr_id3_r <= rcsr_id2_r; // @[memory.scala 359:21]
    end
    if (reset) begin // @[memory.scala 340:30]
      special3_r <= 2'h0; // @[memory.scala 340:30]
    end else if (hs2) begin // @[memory.scala 349:14]
      special3_r <= special2_r; // @[memory.scala 360:21]
    end
    if (reset) begin // @[memory.scala 341:30]
      is_mmio_r <= 1'h0; // @[memory.scala 341:30]
    end else if (hs2) begin // @[memory.scala 349:14]
      is_mmio_r <= is_dc_r & paddr2_r < 32'h80000000; // @[memory.scala 362:21]
    end
    if (reset) begin // @[memory.scala 342:30]
      recov3_r <= 1'h0; // @[memory.scala 342:30]
    end else if (hs2) begin // @[memory.scala 349:14]
      recov3_r <= recov2_r; // @[memory.scala 361:21]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  drop2_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  stall2_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  inst1_r = _RAND_2[31:0];
  _RAND_3 = {2{`RANDOM}};
  pc1_r = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  excep1_r_cause = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  excep1_r_tval = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  excep1_r_en = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  excep1_r_pc = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  excep1_r_etype = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  ctrl1_r_dcMode = _RAND_9[4:0];
  _RAND_10 = {2{`RANDOM}};
  mem_addr1_r = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mem_data1_r = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  dst1_r = _RAND_12[4:0];
  _RAND_13 = {2{`RANDOM}};
  dst_d1_r = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  dst_en1_r = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  csr_id1_r = _RAND_15[11:0];
  _RAND_16 = {2{`RANDOM}};
  csr_d1_r = _RAND_16[63:0];
  _RAND_17 = {1{`RANDOM}};
  csr_en1_r = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  rcsr_id1_r = _RAND_18[11:0];
  _RAND_19 = {1{`RANDOM}};
  special1_r = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  indi1_r = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  recov1_r = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid1_r = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  is_tlb_r = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  drop_tlb = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid2_r = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid3_r = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  ctrl2_r_dcMode = _RAND_27[4:0];
  _RAND_28 = {1{`RANDOM}};
  drop_dc = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  inst2_r = _RAND_29[31:0];
  _RAND_30 = {2{`RANDOM}};
  pc2_r = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  excep2_r_cause = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  excep2_r_tval = _RAND_32[63:0];
  _RAND_33 = {1{`RANDOM}};
  excep2_r_en = _RAND_33[0:0];
  _RAND_34 = {2{`RANDOM}};
  excep2_r_pc = _RAND_34[63:0];
  _RAND_35 = {1{`RANDOM}};
  excep2_r_etype = _RAND_35[1:0];
  _RAND_36 = {2{`RANDOM}};
  mem_data2_r = _RAND_36[63:0];
  _RAND_37 = {1{`RANDOM}};
  dst2_r = _RAND_37[4:0];
  _RAND_38 = {2{`RANDOM}};
  dst_d2_r = _RAND_38[63:0];
  _RAND_39 = {1{`RANDOM}};
  dst_en2_r = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  csr_id2_r = _RAND_40[11:0];
  _RAND_41 = {2{`RANDOM}};
  csr_d2_r = _RAND_41[63:0];
  _RAND_42 = {1{`RANDOM}};
  csr_en2_r = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  rcsr_id2_r = _RAND_43[11:0];
  _RAND_44 = {1{`RANDOM}};
  special2_r = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  paddr2_r = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  recov2_r = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  dc_hs_r = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  lr_addr_r = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  lr_valid_r = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  inst3_r = _RAND_50[31:0];
  _RAND_51 = {2{`RANDOM}};
  pc3_r = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  excep3_r_cause = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  excep3_r_tval = _RAND_53[63:0];
  _RAND_54 = {1{`RANDOM}};
  excep3_r_en = _RAND_54[0:0];
  _RAND_55 = {2{`RANDOM}};
  excep3_r_pc = _RAND_55[63:0];
  _RAND_56 = {1{`RANDOM}};
  excep3_r_etype = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  dst3_r = _RAND_57[4:0];
  _RAND_58 = {2{`RANDOM}};
  dst_d3_r = _RAND_58[63:0];
  _RAND_59 = {1{`RANDOM}};
  dst_en3_r = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  csr_id3_r = _RAND_60[11:0];
  _RAND_61 = {2{`RANDOM}};
  csr_d3_r = _RAND_61[63:0];
  _RAND_62 = {1{`RANDOM}};
  csr_en3_r = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  rcsr_id3_r = _RAND_63[11:0];
  _RAND_64 = {1{`RANDOM}};
  special3_r = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  is_mmio_r = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  recov3_r = _RAND_66[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_Writeback(
  input         clock,
  input         reset,
  input  [31:0] io_mem2rb_inst,
  input  [63:0] io_mem2rb_pc,
  input  [63:0] io_mem2rb_excep_cause,
  input  [63:0] io_mem2rb_excep_tval,
  input         io_mem2rb_excep_en,
  input  [63:0] io_mem2rb_excep_pc,
  input  [1:0]  io_mem2rb_excep_etype,
  input  [11:0] io_mem2rb_csr_id,
  input  [63:0] io_mem2rb_csr_d,
  input         io_mem2rb_csr_en,
  input  [4:0]  io_mem2rb_dst,
  input  [63:0] io_mem2rb_dst_d,
  input         io_mem2rb_dst_en,
  input  [11:0] io_mem2rb_rcsr_id,
  input  [1:0]  io_mem2rb_special,
  input         io_mem2rb_is_mmio,
  output        io_mem2rb_drop,
  output        io_mem2rb_stall,
  input         io_mem2rb_recov,
  input         io_mem2rb_valid,
  output        io_mem2rb_ready,
  output [4:0]  io_wReg_id,
  output [63:0] io_wReg_data,
  output        io_wReg_en,
  output [11:0] io_wCsr_id,
  output [63:0] io_wCsr_data,
  output        io_wCsr_en,
  output [63:0] io_excep_cause,
  output [63:0] io_excep_tval,
  output        io_excep_en,
  output [63:0] io_excep_pc,
  output [1:0]  io_excep_etype,
  output [63:0] io_wb2if_seq_pc,
  output        io_wb2if_valid,
  output        io_recov,
  output        io_flush_tlb,
  output        io_flush_cache
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  recov_r; // @[writeback.scala 22:30]
  reg [63:0] forceJmp_seq_pc; // @[writeback.scala 25:30]
  reg  forceJmp_valid; // @[writeback.scala 25:30]
  reg  tlb_r; // @[writeback.scala 26:30]
  reg  cache_r; // @[writeback.scala 27:30]
  wire  _T_4 = io_mem2rb_special != 2'h0 | io_mem2rb_recov & ~io_mem2rb_excep_en; // @[writeback.scala 67:44]
  wire [63:0] _forceJmp_seq_pc_T_1 = io_mem2rb_pc + 64'h4; // @[writeback.scala 69:49]
  wire  _T_5 = io_mem2rb_special == 2'h1; // @[writeback.scala 70:40]
  wire  _T_6 = io_mem2rb_special == 2'h2; // @[writeback.scala 72:46]
  wire  _GEN_2 = io_mem2rb_special == 2'h1 ? 1'h0 : _T_6; // @[writeback.scala 70:60 writeback.scala 32:21]
  wire  _GEN_5 = (io_mem2rb_special != 2'h0 | io_mem2rb_recov & ~io_mem2rb_excep_en) & _T_5; // @[writeback.scala 67:88 writeback.scala 33:21]
  wire  _GEN_6 = (io_mem2rb_special != 2'h0 | io_mem2rb_recov & ~io_mem2rb_excep_en) & _GEN_2; // @[writeback.scala 67:88 writeback.scala 32:21]
  wire  _GEN_13 = io_mem2rb_valid & io_mem2rb_recov; // @[writeback.scala 56:30 writeback.scala 64:21 writeback.scala 24:32]
  wire  _GEN_19 = io_mem2rb_valid & _T_4; // @[writeback.scala 56:30 writeback.scala 34:21]
  wire  _GEN_21 = io_mem2rb_valid & _GEN_5; // @[writeback.scala 56:30 writeback.scala 33:21]
  wire  _GEN_22 = io_mem2rb_valid & _GEN_6; // @[writeback.scala 56:30 writeback.scala 32:21]
  assign io_mem2rb_drop = 1'h0; // @[writeback.scala 38:21]
  assign io_mem2rb_stall = 1'h0; // @[writeback.scala 54:21]
  assign io_mem2rb_ready = io_mem2rb_valid; // @[writeback.scala 55:18 writeback.scala 53:21]
  assign io_wReg_id = io_mem2rb_dst; // @[writeback.scala 42:21]
  assign io_wReg_data = io_mem2rb_dst_d; // @[writeback.scala 43:21]
  assign io_wReg_en = io_mem2rb_valid & io_mem2rb_dst_en; // @[writeback.scala 56:30 writeback.scala 58:29 writeback.scala 44:21]
  assign io_wCsr_id = io_mem2rb_csr_id; // @[writeback.scala 45:21]
  assign io_wCsr_data = io_mem2rb_csr_d; // @[writeback.scala 46:21]
  assign io_wCsr_en = io_mem2rb_valid & io_mem2rb_csr_en; // @[writeback.scala 56:30 writeback.scala 59:29 writeback.scala 47:21]
  assign io_excep_cause = io_mem2rb_excep_cause; // @[writeback.scala 48:21]
  assign io_excep_tval = io_mem2rb_excep_tval; // @[writeback.scala 48:21]
  assign io_excep_en = io_mem2rb_valid & io_mem2rb_excep_en; // @[writeback.scala 56:30 writeback.scala 60:29 writeback.scala 49:21]
  assign io_excep_pc = io_mem2rb_excep_pc; // @[writeback.scala 48:21]
  assign io_excep_etype = io_mem2rb_excep_etype; // @[writeback.scala 48:21]
  assign io_wb2if_seq_pc = forceJmp_seq_pc; // @[writeback.scala 52:21]
  assign io_wb2if_valid = forceJmp_valid; // @[writeback.scala 52:21]
  assign io_recov = recov_r; // @[writeback.scala 39:21]
  assign io_flush_tlb = tlb_r; // @[writeback.scala 50:21]
  assign io_flush_cache = cache_r; // @[writeback.scala 51:21]
  always @(posedge clock) begin
    if (reset) begin // @[writeback.scala 22:30]
      recov_r <= 1'h0; // @[writeback.scala 22:30]
    end else begin
      recov_r <= _GEN_13;
    end
    if (reset) begin // @[writeback.scala 25:30]
      forceJmp_seq_pc <= 64'h0; // @[writeback.scala 25:30]
    end else if (io_mem2rb_valid) begin // @[writeback.scala 56:30]
      if (io_mem2rb_special != 2'h0 | io_mem2rb_recov & ~io_mem2rb_excep_en) begin // @[writeback.scala 67:88]
        forceJmp_seq_pc <= _forceJmp_seq_pc_T_1; // @[writeback.scala 69:33]
      end
    end
    if (reset) begin // @[writeback.scala 25:30]
      forceJmp_valid <= 1'h0; // @[writeback.scala 25:30]
    end else begin
      forceJmp_valid <= _GEN_19;
    end
    if (reset) begin // @[writeback.scala 26:30]
      tlb_r <= 1'h0; // @[writeback.scala 26:30]
    end else begin
      tlb_r <= _GEN_22;
    end
    if (reset) begin // @[writeback.scala 27:30]
      cache_r <= 1'h0; // @[writeback.scala 27:30]
    end else begin
      cache_r <= _GEN_21;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  recov_r = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  forceJmp_seq_pc = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  forceJmp_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  tlb_r = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  cache_r = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_Regs(
  input         clock,
  input         reset,
  input  [4:0]  io_rs1_id,
  output [63:0] io_rs1_data,
  input  [4:0]  io_rs2_id,
  output [63:0] io_rs2_data,
  input  [4:0]  io_dst_id,
  input  [63:0] io_dst_data,
  input         io_dst_en
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] regs_0; // @[regs.scala 15:23]
  reg [63:0] regs_1; // @[regs.scala 15:23]
  reg [63:0] regs_2; // @[regs.scala 15:23]
  reg [63:0] regs_3; // @[regs.scala 15:23]
  reg [63:0] regs_4; // @[regs.scala 15:23]
  reg [63:0] regs_5; // @[regs.scala 15:23]
  reg [63:0] regs_6; // @[regs.scala 15:23]
  reg [63:0] regs_7; // @[regs.scala 15:23]
  reg [63:0] regs_8; // @[regs.scala 15:23]
  reg [63:0] regs_9; // @[regs.scala 15:23]
  reg [63:0] regs_10; // @[regs.scala 15:23]
  reg [63:0] regs_11; // @[regs.scala 15:23]
  reg [63:0] regs_12; // @[regs.scala 15:23]
  reg [63:0] regs_13; // @[regs.scala 15:23]
  reg [63:0] regs_14; // @[regs.scala 15:23]
  reg [63:0] regs_15; // @[regs.scala 15:23]
  reg [63:0] regs_16; // @[regs.scala 15:23]
  reg [63:0] regs_17; // @[regs.scala 15:23]
  reg [63:0] regs_18; // @[regs.scala 15:23]
  reg [63:0] regs_19; // @[regs.scala 15:23]
  reg [63:0] regs_20; // @[regs.scala 15:23]
  reg [63:0] regs_21; // @[regs.scala 15:23]
  reg [63:0] regs_22; // @[regs.scala 15:23]
  reg [63:0] regs_23; // @[regs.scala 15:23]
  reg [63:0] regs_24; // @[regs.scala 15:23]
  reg [63:0] regs_25; // @[regs.scala 15:23]
  reg [63:0] regs_26; // @[regs.scala 15:23]
  reg [63:0] regs_27; // @[regs.scala 15:23]
  reg [63:0] regs_28; // @[regs.scala 15:23]
  reg [63:0] regs_29; // @[regs.scala 15:23]
  reg [63:0] regs_30; // @[regs.scala 15:23]
  reg [63:0] regs_31; // @[regs.scala 15:23]
  wire [63:0] _GEN_1 = 5'h1 == io_rs1_id ? regs_1 : regs_0; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_2 = 5'h2 == io_rs1_id ? regs_2 : _GEN_1; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_3 = 5'h3 == io_rs1_id ? regs_3 : _GEN_2; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_4 = 5'h4 == io_rs1_id ? regs_4 : _GEN_3; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_5 = 5'h5 == io_rs1_id ? regs_5 : _GEN_4; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_6 = 5'h6 == io_rs1_id ? regs_6 : _GEN_5; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_7 = 5'h7 == io_rs1_id ? regs_7 : _GEN_6; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_8 = 5'h8 == io_rs1_id ? regs_8 : _GEN_7; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_9 = 5'h9 == io_rs1_id ? regs_9 : _GEN_8; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_10 = 5'ha == io_rs1_id ? regs_10 : _GEN_9; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_11 = 5'hb == io_rs1_id ? regs_11 : _GEN_10; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_12 = 5'hc == io_rs1_id ? regs_12 : _GEN_11; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_13 = 5'hd == io_rs1_id ? regs_13 : _GEN_12; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_14 = 5'he == io_rs1_id ? regs_14 : _GEN_13; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_15 = 5'hf == io_rs1_id ? regs_15 : _GEN_14; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_16 = 5'h10 == io_rs1_id ? regs_16 : _GEN_15; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_17 = 5'h11 == io_rs1_id ? regs_17 : _GEN_16; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_18 = 5'h12 == io_rs1_id ? regs_18 : _GEN_17; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_19 = 5'h13 == io_rs1_id ? regs_19 : _GEN_18; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_20 = 5'h14 == io_rs1_id ? regs_20 : _GEN_19; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_21 = 5'h15 == io_rs1_id ? regs_21 : _GEN_20; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_22 = 5'h16 == io_rs1_id ? regs_22 : _GEN_21; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_23 = 5'h17 == io_rs1_id ? regs_23 : _GEN_22; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_24 = 5'h18 == io_rs1_id ? regs_24 : _GEN_23; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_25 = 5'h19 == io_rs1_id ? regs_25 : _GEN_24; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_26 = 5'h1a == io_rs1_id ? regs_26 : _GEN_25; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_27 = 5'h1b == io_rs1_id ? regs_27 : _GEN_26; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_28 = 5'h1c == io_rs1_id ? regs_28 : _GEN_27; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_29 = 5'h1d == io_rs1_id ? regs_29 : _GEN_28; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_30 = 5'h1e == io_rs1_id ? regs_30 : _GEN_29; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_31 = 5'h1f == io_rs1_id ? regs_31 : _GEN_30; // @[regs.scala 17:23 regs.scala 17:23]
  wire [63:0] _GEN_33 = 5'h1 == io_rs2_id ? regs_1 : regs_0; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_34 = 5'h2 == io_rs2_id ? regs_2 : _GEN_33; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_35 = 5'h3 == io_rs2_id ? regs_3 : _GEN_34; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_36 = 5'h4 == io_rs2_id ? regs_4 : _GEN_35; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_37 = 5'h5 == io_rs2_id ? regs_5 : _GEN_36; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_38 = 5'h6 == io_rs2_id ? regs_6 : _GEN_37; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_39 = 5'h7 == io_rs2_id ? regs_7 : _GEN_38; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_40 = 5'h8 == io_rs2_id ? regs_8 : _GEN_39; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_41 = 5'h9 == io_rs2_id ? regs_9 : _GEN_40; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_42 = 5'ha == io_rs2_id ? regs_10 : _GEN_41; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_43 = 5'hb == io_rs2_id ? regs_11 : _GEN_42; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_44 = 5'hc == io_rs2_id ? regs_12 : _GEN_43; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_45 = 5'hd == io_rs2_id ? regs_13 : _GEN_44; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_46 = 5'he == io_rs2_id ? regs_14 : _GEN_45; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_47 = 5'hf == io_rs2_id ? regs_15 : _GEN_46; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_48 = 5'h10 == io_rs2_id ? regs_16 : _GEN_47; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_49 = 5'h11 == io_rs2_id ? regs_17 : _GEN_48; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_50 = 5'h12 == io_rs2_id ? regs_18 : _GEN_49; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_51 = 5'h13 == io_rs2_id ? regs_19 : _GEN_50; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_52 = 5'h14 == io_rs2_id ? regs_20 : _GEN_51; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_53 = 5'h15 == io_rs2_id ? regs_21 : _GEN_52; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_54 = 5'h16 == io_rs2_id ? regs_22 : _GEN_53; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_55 = 5'h17 == io_rs2_id ? regs_23 : _GEN_54; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_56 = 5'h18 == io_rs2_id ? regs_24 : _GEN_55; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_57 = 5'h19 == io_rs2_id ? regs_25 : _GEN_56; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_58 = 5'h1a == io_rs2_id ? regs_26 : _GEN_57; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_59 = 5'h1b == io_rs2_id ? regs_27 : _GEN_58; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_60 = 5'h1c == io_rs2_id ? regs_28 : _GEN_59; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_61 = 5'h1d == io_rs2_id ? regs_29 : _GEN_60; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_62 = 5'h1e == io_rs2_id ? regs_30 : _GEN_61; // @[regs.scala 18:23 regs.scala 18:23]
  wire [63:0] _GEN_63 = 5'h1f == io_rs2_id ? regs_31 : _GEN_62; // @[regs.scala 18:23 regs.scala 18:23]
  assign io_rs1_data = io_rs1_id == 5'h0 ? 64'h0 : _GEN_31; // @[regs.scala 17:23]
  assign io_rs2_data = io_rs2_id == 5'h0 ? 64'h0 : _GEN_63; // @[regs.scala 18:23]
  always @(posedge clock) begin
    if (reset) begin // @[regs.scala 15:23]
      regs_0 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h0 == io_dst_id) begin // @[regs.scala 20:25]
        regs_0 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_1 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h1 == io_dst_id) begin // @[regs.scala 20:25]
        regs_1 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_2 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h2 == io_dst_id) begin // @[regs.scala 20:25]
        regs_2 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_3 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h3 == io_dst_id) begin // @[regs.scala 20:25]
        regs_3 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_4 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h4 == io_dst_id) begin // @[regs.scala 20:25]
        regs_4 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_5 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h5 == io_dst_id) begin // @[regs.scala 20:25]
        regs_5 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_6 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h6 == io_dst_id) begin // @[regs.scala 20:25]
        regs_6 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_7 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h7 == io_dst_id) begin // @[regs.scala 20:25]
        regs_7 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_8 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h8 == io_dst_id) begin // @[regs.scala 20:25]
        regs_8 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_9 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h9 == io_dst_id) begin // @[regs.scala 20:25]
        regs_9 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_10 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'ha == io_dst_id) begin // @[regs.scala 20:25]
        regs_10 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_11 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'hb == io_dst_id) begin // @[regs.scala 20:25]
        regs_11 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_12 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'hc == io_dst_id) begin // @[regs.scala 20:25]
        regs_12 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_13 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'hd == io_dst_id) begin // @[regs.scala 20:25]
        regs_13 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_14 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'he == io_dst_id) begin // @[regs.scala 20:25]
        regs_14 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_15 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'hf == io_dst_id) begin // @[regs.scala 20:25]
        regs_15 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_16 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h10 == io_dst_id) begin // @[regs.scala 20:25]
        regs_16 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_17 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h11 == io_dst_id) begin // @[regs.scala 20:25]
        regs_17 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_18 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h12 == io_dst_id) begin // @[regs.scala 20:25]
        regs_18 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_19 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h13 == io_dst_id) begin // @[regs.scala 20:25]
        regs_19 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_20 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h14 == io_dst_id) begin // @[regs.scala 20:25]
        regs_20 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_21 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h15 == io_dst_id) begin // @[regs.scala 20:25]
        regs_21 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_22 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h16 == io_dst_id) begin // @[regs.scala 20:25]
        regs_22 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_23 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h17 == io_dst_id) begin // @[regs.scala 20:25]
        regs_23 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_24 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h18 == io_dst_id) begin // @[regs.scala 20:25]
        regs_24 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_25 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h19 == io_dst_id) begin // @[regs.scala 20:25]
        regs_25 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_26 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h1a == io_dst_id) begin // @[regs.scala 20:25]
        regs_26 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_27 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h1b == io_dst_id) begin // @[regs.scala 20:25]
        regs_27 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_28 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h1c == io_dst_id) begin // @[regs.scala 20:25]
        regs_28 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_29 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h1d == io_dst_id) begin // @[regs.scala 20:25]
        regs_29 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_30 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h1e == io_dst_id) begin // @[regs.scala 20:25]
        regs_30 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
    if (reset) begin // @[regs.scala 15:23]
      regs_31 <= 64'h0; // @[regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[regs.scala 19:41]
      if (5'h1f == io_dst_id) begin // @[regs.scala 20:25]
        regs_31 <= io_dst_data; // @[regs.scala 20:25]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regs_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regs_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  regs_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  regs_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  regs_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  regs_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  regs_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  regs_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  regs_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  regs_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  regs_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  regs_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  regs_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  regs_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  regs_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  regs_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  regs_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  regs_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  regs_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  regs_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  regs_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  regs_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  regs_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  regs_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  regs_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  regs_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  regs_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  regs_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  regs_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  regs_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  regs_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  regs_31 = _RAND_31[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_Csrs(
  input         clock,
  input         reset,
  input  [11:0] io_rs_id,
  output [63:0] io_rs_data,
  output        io_rs_is_err,
  input  [11:0] io_rd_id,
  input  [63:0] io_rd_data,
  input         io_rd_en,
  input  [63:0] io_excep_cause,
  input  [63:0] io_excep_tval,
  input         io_excep_en,
  input  [63:0] io_excep_pc,
  input  [1:0]  io_excep_etype,
  output [1:0]  io_mmuState_priv,
  output [63:0] io_mmuState_mstatus,
  output [63:0] io_mmuState_satp,
  output [1:0]  io_idState_priv,
  output [63:0] io_reg2if_seq_pc,
  output        io_reg2if_valid,
  output        io_intr_out_en,
  output [63:0] io_intr_out_cause,
  input         io_clint_raise,
  input         io_clint_clear,
  input         io_plic_m_raise,
  input         io_plic_m_clear,
  input         io_plic_s_raise,
  input         io_plic_s_clear,
  output [63:0] io_updateNextPc_seq_pc,
  output        io_updateNextPc_valid,
  input         io_intr_msip_raise,
  input         io_intr_msip_clear
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] priv; // @[regs.scala 42:30]
  reg [63:0] misa; // @[regs.scala 43:30]
  reg [63:0] mstatus; // @[regs.scala 44:30]
  reg [63:0] mepc; // @[regs.scala 45:30]
  reg [63:0] mtval; // @[regs.scala 46:30]
  reg [63:0] mscratch; // @[regs.scala 47:30]
  reg [63:0] mcause; // @[regs.scala 48:30]
  reg [63:0] mtvec; // @[regs.scala 49:30]
  reg [63:0] mie; // @[regs.scala 50:30]
  reg [63:0] mip; // @[regs.scala 51:30]
  reg [63:0] medeleg; // @[regs.scala 52:30]
  reg [63:0] mideleg; // @[regs.scala 53:30]
  reg [31:0] mcounteren; // @[regs.scala 54:30]
  reg [31:0] scounteren; // @[regs.scala 55:30]
  reg [63:0] sepc; // @[regs.scala 56:30]
  reg [63:0] stval; // @[regs.scala 57:30]
  reg [63:0] sscratch; // @[regs.scala 58:30]
  reg [63:0] stvec; // @[regs.scala 59:30]
  reg [63:0] satp; // @[regs.scala 60:30]
  reg [63:0] scause; // @[regs.scala 61:30]
  reg [63:0] pmpaddr0; // @[regs.scala 62:30]
  reg [63:0] pmpaddr1; // @[regs.scala 63:30]
  reg [63:0] pmpaddr2; // @[regs.scala 64:30]
  reg [63:0] pmpaddr3; // @[regs.scala 65:30]
  reg [63:0] uscratch; // @[regs.scala 66:30]
  reg [63:0] mhartid; // @[regs.scala 68:30]
  wire [63:0] sstatus = mstatus & 64'h80000003000de122; // @[regs.scala 69:31]
  reg [63:0] forceJmp_seq_pc; // @[regs.scala 75:34]
  reg  forceJmp_valid; // @[regs.scala 75:34]
  wire  priv_lo = sstatus[8]; // @[regs.scala 85:48]
  wire [1:0] _priv_T = {1'h0,priv_lo}; // @[Cat.scala 30:58]
  wire [54:0] new_sstatus_hi_hi_hi = sstatus[63:9]; // @[regs.scala 86:37]
  wire [1:0] new_sstatus_hi_lo_hi = sstatus[7:6]; // @[regs.scala 86:57]
  wire [2:0] new_sstatus_lo_hi_hi = sstatus[4:2]; // @[regs.scala 86:76]
  wire  new_sstatus_lo_hi_lo = sstatus[5]; // @[regs.scala 86:85]
  wire  new_sstatus_lo_lo = sstatus[0]; // @[regs.scala 86:92]
  wire [63:0] new_sstatus = {new_sstatus_hi_hi_hi,1'h0,new_sstatus_hi_lo_hi,1'h1,new_sstatus_lo_hi_hi,
    new_sstatus_lo_hi_lo,new_sstatus_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] _mstatus_T_1 = mstatus & 64'hfffffffffff21edd; // @[common.scala 201:17]
  wire [63:0] _mstatus_T_2 = new_sstatus & 64'hde122; // @[common.scala 201:36]
  wire [63:0] _mstatus_T_3 = _mstatus_T_1 | _mstatus_T_2; // @[common.scala 201:26]
  wire [50:0] new_mstatus_hi_hi_hi = mstatus[63:13]; // @[regs.scala 93:37]
  wire [2:0] new_mstatus_hi_lo_hi = mstatus[10:8]; // @[regs.scala 93:55]
  wire [2:0] new_mstatus_lo_hi_hi = mstatus[6:4]; // @[regs.scala 93:75]
  wire  new_mstatus_lo_hi_lo = mstatus[7]; // @[regs.scala 93:84]
  wire [2:0] new_mstatus_lo_lo = mstatus[2:0]; // @[regs.scala 93:91]
  wire [63:0] new_mstatus = {new_mstatus_hi_hi_hi,2'h0,new_mstatus_hi_lo_hi,1'h1,new_mstatus_lo_hi_hi,
    new_mstatus_lo_hi_lo,new_mstatus_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] deleg = io_excep_cause[63] ? mideleg : medeleg; // @[regs.scala 97:28]
  wire  _T_2 = priv <= 2'h1; // @[regs.scala 98:23]
  wire [63:0] _T_4 = deleg >> io_excep_cause[62:0]; // @[regs.scala 98:40]
  wire [65:0] _GEN_550 = {io_excep_cause, 2'h0}; // @[regs.scala 99:66]
  wire [66:0] _seq_pc_T_2 = {{1'd0}, _GEN_550}; // @[regs.scala 99:66]
  wire [66:0] _seq_pc_T_3 = stvec[1] ? _seq_pc_T_2 : 67'h0; // @[regs.scala 99:41]
  wire [66:0] _GEN_551 = {{3'd0}, stvec}; // @[regs.scala 99:36]
  wire [66:0] seq_pc = _GEN_551 + _seq_pc_T_3; // @[regs.scala 99:36]
  wire  new_sstatus_hi_hi_lo = priv[0]; // @[regs.scala 105:53]
  wire  new_sstatus_hi_lo_lo = sstatus[1]; // @[regs.scala 105:69]
  wire [63:0] new_sstatus_1 = {new_sstatus_hi_hi_hi,new_sstatus_hi_hi_lo,new_sstatus_hi_lo_hi,new_sstatus_hi_lo_lo,
    new_sstatus_lo_hi_hi,1'h0,new_sstatus_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] _mstatus_T_6 = new_sstatus_1 & 64'hde122; // @[common.scala 201:36]
  wire [63:0] _mstatus_T_7 = _mstatus_T_1 | _mstatus_T_6; // @[common.scala 201:26]
  wire [66:0] _seq_pc_T_7 = mtvec[1] ? _seq_pc_T_2 : 67'h0; // @[regs.scala 110:46]
  wire [66:0] _GEN_553 = {{3'd0}, mtvec}; // @[regs.scala 110:41]
  wire [66:0] seq_pc_1 = _GEN_553 + _seq_pc_T_7; // @[regs.scala 110:41]
  wire  new_mstatus_hi_lo_lo = mstatus[3]; // @[regs.scala 116:73]
  wire [63:0] new_mstatus_1 = {new_mstatus_hi_hi_hi,priv,new_mstatus_hi_lo_hi,new_mstatus_hi_lo_lo,new_mstatus_lo_hi_hi,1'h0
    ,new_mstatus_lo_lo}; // @[Cat.scala 30:58]
  wire [66:0] _GEN_0 = priv <= 2'h1 & _T_4[0] ? seq_pc : seq_pc_1; // @[regs.scala 98:54 regs.scala 100:33 regs.scala 111:33]
  wire [63:0] _GEN_2 = priv <= 2'h1 & _T_4[0] ? io_excep_cause : scause; // @[regs.scala 98:54 regs.scala 102:33 regs.scala 61:30]
  wire [63:0] _GEN_3 = priv <= 2'h1 & _T_4[0] ? io_excep_pc : sepc; // @[regs.scala 98:54 regs.scala 103:33 regs.scala 56:30]
  wire [63:0] _GEN_4 = priv <= 2'h1 & _T_4[0] ? _mstatus_T_7 : new_mstatus_1; // @[regs.scala 98:54 regs.scala 106:33 regs.scala 117:33]
  wire [63:0] _GEN_5 = priv <= 2'h1 & _T_4[0] ? io_excep_tval : stval; // @[regs.scala 98:54 regs.scala 107:33 regs.scala 57:30]
  wire [1:0] _GEN_6 = priv <= 2'h1 & _T_4[0] ? 2'h1 : 2'h3; // @[regs.scala 98:54 regs.scala 108:33 regs.scala 119:33]
  wire [63:0] _GEN_7 = priv <= 2'h1 & _T_4[0] ? mcause : io_excep_cause; // @[regs.scala 98:54 regs.scala 48:30 regs.scala 113:33]
  wire [63:0] _GEN_8 = priv <= 2'h1 & _T_4[0] ? mepc : io_excep_pc; // @[regs.scala 98:54 regs.scala 45:30 regs.scala 114:33]
  wire [63:0] _GEN_9 = priv <= 2'h1 & _T_4[0] ? mtval : io_excep_tval; // @[regs.scala 98:54 regs.scala 46:30 regs.scala 118:33]
  wire [66:0] _GEN_10 = io_excep_etype == 2'h3 ? {{3'd0}, mepc} : _GEN_0; // @[regs.scala 88:50 regs.scala 89:29]
  wire [63:0] _GEN_13 = io_excep_etype == 2'h3 ? new_mstatus : _GEN_4; // @[regs.scala 88:50 regs.scala 94:29]
  wire [63:0] _GEN_14 = io_excep_etype == 2'h3 ? scause : _GEN_2; // @[regs.scala 88:50 regs.scala 61:30]
  wire [63:0] _GEN_15 = io_excep_etype == 2'h3 ? sepc : _GEN_3; // @[regs.scala 88:50 regs.scala 56:30]
  wire [63:0] _GEN_16 = io_excep_etype == 2'h3 ? stval : _GEN_5; // @[regs.scala 88:50 regs.scala 57:30]
  wire [63:0] _GEN_17 = io_excep_etype == 2'h3 ? mcause : _GEN_7; // @[regs.scala 88:50 regs.scala 48:30]
  wire [63:0] _GEN_18 = io_excep_etype == 2'h3 ? mepc : _GEN_8; // @[regs.scala 88:50 regs.scala 45:30]
  wire [63:0] _GEN_19 = io_excep_etype == 2'h3 ? mtval : _GEN_9; // @[regs.scala 88:50 regs.scala 46:30]
  wire [66:0] _GEN_20 = io_excep_etype == 2'h2 ? {{3'd0}, sepc} : _GEN_10; // @[regs.scala 81:44 regs.scala 82:29]
  wire [63:0] _GEN_23 = io_excep_etype == 2'h2 ? _mstatus_T_3 : _GEN_13; // @[regs.scala 81:44 regs.scala 87:29]
  wire [63:0] _GEN_24 = io_excep_etype == 2'h2 ? scause : _GEN_14; // @[regs.scala 81:44 regs.scala 61:30]
  wire [63:0] _GEN_25 = io_excep_etype == 2'h2 ? sepc : _GEN_15; // @[regs.scala 81:44 regs.scala 56:30]
  wire [63:0] _GEN_26 = io_excep_etype == 2'h2 ? stval : _GEN_16; // @[regs.scala 81:44 regs.scala 57:30]
  wire [63:0] _GEN_27 = io_excep_etype == 2'h2 ? mcause : _GEN_17; // @[regs.scala 81:44 regs.scala 48:30]
  wire [63:0] _GEN_28 = io_excep_etype == 2'h2 ? mepc : _GEN_18; // @[regs.scala 81:44 regs.scala 45:30]
  wire [63:0] _GEN_29 = io_excep_etype == 2'h2 ? mtval : _GEN_19; // @[regs.scala 81:44 regs.scala 46:30]
  wire [66:0] _GEN_30 = io_excep_en ? _GEN_20 : {{3'd0}, forceJmp_seq_pc}; // @[regs.scala 80:22 regs.scala 75:34]
  wire [63:0] _GEN_33 = io_excep_en ? _GEN_23 : mstatus; // @[regs.scala 80:22 regs.scala 44:30]
  wire [63:0] _GEN_34 = io_excep_en ? _GEN_24 : scause; // @[regs.scala 80:22 regs.scala 61:30]
  wire [63:0] _GEN_35 = io_excep_en ? _GEN_25 : sepc; // @[regs.scala 80:22 regs.scala 56:30]
  wire [63:0] _GEN_36 = io_excep_en ? _GEN_26 : stval; // @[regs.scala 80:22 regs.scala 57:30]
  wire [63:0] _GEN_37 = io_excep_en ? _GEN_27 : mcause; // @[regs.scala 80:22 regs.scala 48:30]
  wire [63:0] _GEN_38 = io_excep_en ? _GEN_28 : mepc; // @[regs.scala 80:22 regs.scala 45:30]
  wire [63:0] _GEN_39 = io_excep_en ? _GEN_29 : mtval; // @[regs.scala 80:22 regs.scala 46:30]
  reg  intr_out_r_en; // @[regs.scala 124:29]
  reg [63:0] intr_out_r_cause; // @[regs.scala 124:29]
  reg  intr_seip; // @[regs.scala 126:28]
  wire [63:0] _mip_T_2 = mip & 64'hffffffffffffff7f; // @[common.scala 201:17]
  wire [63:0] _mip_T_4 = _mip_T_2 | 64'h80; // @[common.scala 201:26]
  wire [63:0] _GEN_40 = io_clint_raise ? _mip_T_4 : mip; // @[regs.scala 127:25 regs.scala 128:13 regs.scala 51:30]
  wire [63:0] _GEN_41 = io_clint_clear ? _mip_T_2 : _GEN_40; // @[regs.scala 130:25 regs.scala 131:13]
  wire [63:0] _mip_T_11 = mip & 64'hfffffffffffff7ff; // @[common.scala 201:17]
  wire [63:0] _mip_T_13 = _mip_T_11 | 64'h800; // @[common.scala 201:26]
  wire [63:0] _GEN_42 = io_plic_m_raise ? _mip_T_13 : _GEN_41; // @[regs.scala 133:26 regs.scala 134:13]
  wire [63:0] _GEN_43 = io_plic_m_clear ? _mip_T_11 : _GEN_42; // @[regs.scala 136:26 regs.scala 137:13]
  wire  _GEN_44 = io_plic_s_raise | intr_seip; // @[regs.scala 139:26 regs.scala 140:19 regs.scala 126:28]
  wire [63:0] _mip_T_20 = mip & 64'hfffffffffffffff7; // @[common.scala 201:17]
  wire [63:0] _mip_T_22 = _mip_T_20 | 64'h8; // @[common.scala 201:26]
  wire [63:0] _GEN_46 = io_intr_msip_raise ? _mip_T_22 : _GEN_43; // @[regs.scala 145:29 regs.scala 146:13]
  wire [63:0] _GEN_47 = io_intr_msip_clear ? _mip_T_20 : _GEN_46; // @[regs.scala 148:29 regs.scala 149:13]
  wire [9:0] _GEN_554 = {intr_seip, 9'h0}; // @[regs.scala 151:42]
  wire [15:0] _pending_int_T = {{6'd0}, _GEN_554}; // @[regs.scala 151:42]
  wire [63:0] _GEN_555 = {{48'd0}, _pending_int_T}; // @[regs.scala 151:29]
  wire [63:0] _pending_int_T_1 = mip | _GEN_555; // @[regs.scala 151:29]
  wire [63:0] pending_int = _pending_int_T_1 & mie; // @[regs.scala 151:59]
  wire  m_enable = priv < 2'h3 | priv == 2'h3 & new_mstatus_hi_lo_lo; // @[regs.scala 152:35]
  wire [63:0] _enable_int_m_T = ~mideleg; // @[regs.scala 153:38]
  wire [63:0] _enable_int_m_T_1 = pending_int & _enable_int_m_T; // @[regs.scala 153:36]
  wire [63:0] _enable_int_m_T_4 = m_enable ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] enable_int_m = _enable_int_m_T_1 & _enable_int_m_T_4; // @[regs.scala 153:47]
  wire  s_enable = _T_2 & mstatus[1]; // @[regs.scala 154:36]
  wire [63:0] _enable_int_s_T = pending_int & mideleg; // @[regs.scala 155:36]
  wire [63:0] _enable_int_s_T_3 = s_enable ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] enable_int_s = _enable_int_s_T & _enable_int_s_T_3; // @[regs.scala 155:46]
  wire [63:0] enable_int = enable_int_m != 64'h0 ? enable_int_m : enable_int_s; // @[regs.scala 156:25]
  wire [5:0] _intr_out_r_cause_T_6 = enable_int[5] ? 6'h5 : 6'h3f; // @[Mux.scala 47:69]
  wire [5:0] _intr_out_r_cause_T_7 = enable_int[1] ? 6'h1 : _intr_out_r_cause_T_6; // @[Mux.scala 47:69]
  wire [5:0] _intr_out_r_cause_T_8 = enable_int[9] ? 6'h9 : _intr_out_r_cause_T_7; // @[Mux.scala 47:69]
  wire [5:0] _intr_out_r_cause_T_9 = enable_int[7] ? 6'h7 : _intr_out_r_cause_T_8; // @[Mux.scala 47:69]
  wire [5:0] _intr_out_r_cause_T_10 = enable_int[3] ? 6'h3 : _intr_out_r_cause_T_9; // @[Mux.scala 47:69]
  wire [5:0] _intr_out_r_cause_T_11 = enable_int[11] ? 6'hb : _intr_out_r_cause_T_10; // @[Mux.scala 47:69]
  wire [63:0] _GEN_556 = {{58'd0}, _intr_out_r_cause_T_11}; // @[regs.scala 168:8]
  wire [63:0] _intr_out_r_cause_T_13 = _GEN_556 | 64'h8000000000000000; // @[regs.scala 168:8]
  wire [63:0] _io_rs_data_T = mie & mideleg; // @[regs.scala 212:27]
  wire [63:0] _io_rs_data_T_1 = mip & 64'h222; // @[regs.scala 214:27]
  wire [63:0] _GEN_48 = io_rs_id == 12'hf14 ? mhartid : 64'h0; // @[regs.scala 227:41 regs.scala 228:20 regs.scala 230:25]
  wire  _GEN_49 = io_rs_id == 12'hf14 ? 1'h0 : 1'h1; // @[regs.scala 227:41 regs.scala 170:21 regs.scala 231:25]
  wire [63:0] _GEN_50 = io_rs_id == 12'h40 ? uscratch : _GEN_48; // @[regs.scala 225:42 regs.scala 226:20]
  wire  _GEN_51 = io_rs_id == 12'h40 ? 1'h0 : _GEN_49; // @[regs.scala 225:42 regs.scala 170:21]
  wire [63:0] _GEN_52 = io_rs_id == 12'h3a0 ? pmpaddr3 : _GEN_50; // @[regs.scala 223:41 regs.scala 224:20]
  wire  _GEN_53 = io_rs_id == 12'h3a0 ? 1'h0 : _GEN_51; // @[regs.scala 223:41 regs.scala 170:21]
  wire [63:0] _GEN_54 = io_rs_id == 12'h3b3 ? pmpaddr3 : _GEN_52; // @[regs.scala 221:42 regs.scala 222:20]
  wire  _GEN_55 = io_rs_id == 12'h3b3 ? 1'h0 : _GEN_53; // @[regs.scala 221:42 regs.scala 170:21]
  wire [63:0] _GEN_56 = io_rs_id == 12'h3b2 ? pmpaddr2 : _GEN_54; // @[regs.scala 219:42 regs.scala 220:20]
  wire  _GEN_57 = io_rs_id == 12'h3b2 ? 1'h0 : _GEN_55; // @[regs.scala 219:42 regs.scala 170:21]
  wire [63:0] _GEN_58 = io_rs_id == 12'h3b1 ? pmpaddr1 : _GEN_56; // @[regs.scala 217:42 regs.scala 218:20]
  wire  _GEN_59 = io_rs_id == 12'h3b1 ? 1'h0 : _GEN_57; // @[regs.scala 217:42 regs.scala 170:21]
  wire [63:0] _GEN_60 = io_rs_id == 12'h3b0 ? pmpaddr0 : _GEN_58; // @[regs.scala 215:42 regs.scala 216:20]
  wire  _GEN_61 = io_rs_id == 12'h3b0 ? 1'h0 : _GEN_59; // @[regs.scala 215:42 regs.scala 170:21]
  wire [63:0] _GEN_62 = io_rs_id == 12'h144 ? _io_rs_data_T_1 : _GEN_60; // @[regs.scala 213:37 regs.scala 214:20]
  wire  _GEN_63 = io_rs_id == 12'h144 ? 1'h0 : _GEN_61; // @[regs.scala 213:37 regs.scala 170:21]
  wire [63:0] _GEN_64 = io_rs_id == 12'h104 ? _io_rs_data_T : _GEN_62; // @[regs.scala 211:37 regs.scala 212:20]
  wire  _GEN_65 = io_rs_id == 12'h104 ? 1'h0 : _GEN_63; // @[regs.scala 211:37 regs.scala 170:21]
  wire [63:0] _GEN_66 = io_rs_id == 12'h100 ? sstatus : _GEN_64; // @[regs.scala 209:41 regs.scala 210:20]
  wire  _GEN_67 = io_rs_id == 12'h100 ? 1'h0 : _GEN_65; // @[regs.scala 209:41 regs.scala 170:21]
  wire [63:0] _GEN_68 = io_rs_id == 12'h142 ? scause : _GEN_66; // @[regs.scala 207:40 regs.scala 208:20]
  wire  _GEN_69 = io_rs_id == 12'h142 ? 1'h0 : _GEN_67; // @[regs.scala 207:40 regs.scala 170:21]
  wire [63:0] _GEN_70 = io_rs_id == 12'h180 ? satp : _GEN_68; // @[regs.scala 205:38 regs.scala 206:20]
  wire  _GEN_71 = io_rs_id == 12'h180 ? 1'h0 : _GEN_69; // @[regs.scala 205:38 regs.scala 170:21]
  wire [63:0] _GEN_72 = io_rs_id == 12'h105 ? stvec : _GEN_70; // @[regs.scala 203:39 regs.scala 204:20]
  wire  _GEN_73 = io_rs_id == 12'h105 ? 1'h0 : _GEN_71; // @[regs.scala 203:39 regs.scala 170:21]
  wire [63:0] _GEN_74 = io_rs_id == 12'h140 ? sscratch : _GEN_72; // @[regs.scala 201:42 regs.scala 202:20]
  wire  _GEN_75 = io_rs_id == 12'h140 ? 1'h0 : _GEN_73; // @[regs.scala 201:42 regs.scala 170:21]
  wire [63:0] _GEN_76 = io_rs_id == 12'h143 ? stval : _GEN_74; // @[regs.scala 199:39 regs.scala 200:20]
  wire  _GEN_77 = io_rs_id == 12'h143 ? 1'h0 : _GEN_75; // @[regs.scala 199:39 regs.scala 170:21]
  wire [63:0] _GEN_78 = io_rs_id == 12'h141 ? sepc : _GEN_76; // @[regs.scala 197:38 regs.scala 198:20]
  wire  _GEN_79 = io_rs_id == 12'h141 ? 1'h0 : _GEN_77; // @[regs.scala 197:38 regs.scala 170:21]
  wire [63:0] _GEN_80 = io_rs_id == 12'h106 ? {{32'd0}, scounteren} : _GEN_78; // @[regs.scala 195:44 regs.scala 196:20]
  wire  _GEN_81 = io_rs_id == 12'h106 ? 1'h0 : _GEN_79; // @[regs.scala 195:44 regs.scala 170:21]
  wire [63:0] _GEN_82 = io_rs_id == 12'h306 ? {{32'd0}, mcounteren} : _GEN_80; // @[regs.scala 193:44 regs.scala 194:20]
  wire  _GEN_83 = io_rs_id == 12'h306 ? 1'h0 : _GEN_81; // @[regs.scala 193:44 regs.scala 170:21]
  wire [63:0] _GEN_84 = io_rs_id == 12'h303 ? mideleg : _GEN_82; // @[regs.scala 191:41 regs.scala 192:20]
  wire  _GEN_85 = io_rs_id == 12'h303 ? 1'h0 : _GEN_83; // @[regs.scala 191:41 regs.scala 170:21]
  wire [63:0] _GEN_86 = io_rs_id == 12'h302 ? medeleg : _GEN_84; // @[regs.scala 189:41 regs.scala 190:20]
  wire  _GEN_87 = io_rs_id == 12'h302 ? 1'h0 : _GEN_85; // @[regs.scala 189:41 regs.scala 170:21]
  wire [63:0] _GEN_88 = io_rs_id == 12'h342 ? mcause : _GEN_86; // @[regs.scala 187:40 regs.scala 188:20]
  wire  _GEN_89 = io_rs_id == 12'h342 ? 1'h0 : _GEN_87; // @[regs.scala 187:40 regs.scala 170:21]
  wire [63:0] _GEN_90 = io_rs_id == 12'h344 ? mip : _GEN_88; // @[regs.scala 185:37 regs.scala 186:20]
  wire  _GEN_91 = io_rs_id == 12'h344 ? 1'h0 : _GEN_89; // @[regs.scala 185:37 regs.scala 170:21]
  wire [63:0] _GEN_92 = io_rs_id == 12'h304 ? mie : _GEN_90; // @[regs.scala 183:37 regs.scala 184:20]
  wire  _GEN_93 = io_rs_id == 12'h304 ? 1'h0 : _GEN_91; // @[regs.scala 183:37 regs.scala 170:21]
  wire [63:0] _GEN_94 = io_rs_id == 12'h305 ? mtvec : _GEN_92; // @[regs.scala 181:39 regs.scala 182:20]
  wire  _GEN_95 = io_rs_id == 12'h305 ? 1'h0 : _GEN_93; // @[regs.scala 181:39 regs.scala 170:21]
  wire [63:0] _GEN_96 = io_rs_id == 12'h340 ? mscratch : _GEN_94; // @[regs.scala 179:42 regs.scala 180:20]
  wire  _GEN_97 = io_rs_id == 12'h340 ? 1'h0 : _GEN_95; // @[regs.scala 179:42 regs.scala 170:21]
  wire [63:0] _GEN_98 = io_rs_id == 12'h343 ? mtval : _GEN_96; // @[regs.scala 177:39 regs.scala 178:20]
  wire  _GEN_99 = io_rs_id == 12'h343 ? 1'h0 : _GEN_97; // @[regs.scala 177:39 regs.scala 170:21]
  wire [63:0] _GEN_100 = io_rs_id == 12'h341 ? mepc : _GEN_98; // @[regs.scala 175:38 regs.scala 176:20]
  wire  _GEN_101 = io_rs_id == 12'h341 ? 1'h0 : _GEN_99; // @[regs.scala 175:38 regs.scala 170:21]
  wire [63:0] _GEN_102 = io_rs_id == 12'h300 ? mstatus : _GEN_100; // @[regs.scala 173:41 regs.scala 174:20]
  wire  _GEN_103 = io_rs_id == 12'h300 ? 1'h0 : _GEN_101; // @[regs.scala 173:41 regs.scala 170:21]
  wire [63:0] new_mstatus_2 = io_rd_data & 64'h7e7faa; // @[regs.scala 237:38]
  wire [63:0] sd = io_rd_data[14:13] == 2'h3 | io_rd_data[16:15] == 2'h3 ? 64'h8000000000000000 : 64'h0; // @[regs.scala 238:30]
  wire [63:0] _mstatus_T_9 = new_mstatus_2 | sd; // @[regs.scala 239:86]
  wire [63:0] _mstatus_T_11 = mstatus & 64'h7fffffffff818055; // @[common.scala 201:17]
  wire [63:0] _mstatus_T_12 = _mstatus_T_9 & 64'h80000000007e7faa; // @[common.scala 201:36]
  wire [63:0] _mstatus_T_13 = _mstatus_T_11 | _mstatus_T_12; // @[common.scala 201:26]
  wire [63:0] _mip_T_28 = mip & 64'hffffffffffffffdd; // @[common.scala 201:17]
  wire [63:0] _mip_T_29 = io_rd_data & 64'h22; // @[common.scala 201:36]
  wire [63:0] _mip_T_30 = _mip_T_28 | _mip_T_29; // @[common.scala 201:26]
  wire [63:0] _mip_T_32 = _mip_T_30 | _GEN_555; // @[regs.scala 251:61]
  wire [63:0] _medeleg_T = io_rd_data & 64'hb309; // @[regs.scala 255:31]
  wire [63:0] _mideleg_T = io_rd_data & 64'h222; // @[regs.scala 257:31]
  wire [63:0] _satp_T_1 = satp & 64'hffff00000000000; // @[common.scala 201:17]
  wire [63:0] _satp_T_2 = io_rd_data & 64'hf0000fffffffffff; // @[common.scala 201:36]
  wire [63:0] _satp_T_3 = _satp_T_1 | _satp_T_2; // @[common.scala 201:26]
  wire [63:0] _new_mstatus_T_2 = io_rd_data & 64'hde122; // @[common.scala 201:36]
  wire [63:0] new_mstatus_3 = _mstatus_T_1 | _new_mstatus_T_2; // @[common.scala 201:26]
  wire [1:0] mstatus_hi = sd[63:62]; // @[regs.scala 277:26]
  wire [61:0] mstatus_lo = new_mstatus_3[61:0]; // @[regs.scala 277:46]
  wire [63:0] _mstatus_T_14 = {mstatus_hi,mstatus_lo}; // @[Cat.scala 30:58]
  wire [63:0] _mie_T_1 = mie & _enable_int_m_T; // @[common.scala 201:17]
  wire [63:0] _mie_T_2 = io_rd_data & mideleg; // @[common.scala 201:36]
  wire [63:0] _mie_T_3 = _mie_T_1 | _mie_T_2; // @[common.scala 201:26]
  wire [63:0] _mip_T_34 = mip & 64'hfffffffffffffddd; // @[common.scala 201:17]
  wire [63:0] _mip_T_36 = _mip_T_34 | _mideleg_T; // @[common.scala 201:26]
  wire [63:0] _pmpaddr0_T = io_rd_data & 64'h3fffffffffffff; // @[regs.scala 283:32]
  wire [63:0] _GEN_106 = io_rd_id == 12'hf14 ? io_rd_data : mhartid; // @[regs.scala 294:41 regs.scala 295:17 regs.scala 68:30]
  wire [63:0] _GEN_107 = io_rd_id == 12'h40 ? io_rd_data : uscratch; // @[regs.scala 292:42 regs.scala 293:18 regs.scala 66:30]
  wire [63:0] _GEN_108 = io_rd_id == 12'h40 ? mhartid : _GEN_106; // @[regs.scala 292:42 regs.scala 68:30]
  wire [63:0] _GEN_110 = io_rd_id == 12'h3a0 ? uscratch : _GEN_107; // @[regs.scala 290:41 regs.scala 66:30]
  wire [63:0] _GEN_111 = io_rd_id == 12'h3a0 ? mhartid : _GEN_108; // @[regs.scala 290:41 regs.scala 68:30]
  wire [63:0] _GEN_112 = io_rd_id == 12'h3b3 ? _pmpaddr0_T : pmpaddr3; // @[regs.scala 288:42 regs.scala 289:18 regs.scala 65:30]
  wire [63:0] _GEN_114 = io_rd_id == 12'h3b3 ? uscratch : _GEN_110; // @[regs.scala 288:42 regs.scala 66:30]
  wire [63:0] _GEN_115 = io_rd_id == 12'h3b3 ? mhartid : _GEN_111; // @[regs.scala 288:42 regs.scala 68:30]
  wire [63:0] _GEN_116 = io_rd_id == 12'h3b2 ? _pmpaddr0_T : pmpaddr2; // @[regs.scala 286:42 regs.scala 287:18 regs.scala 64:30]
  wire [63:0] _GEN_117 = io_rd_id == 12'h3b2 ? pmpaddr3 : _GEN_112; // @[regs.scala 286:42 regs.scala 65:30]
  wire [63:0] _GEN_119 = io_rd_id == 12'h3b2 ? uscratch : _GEN_114; // @[regs.scala 286:42 regs.scala 66:30]
  wire [63:0] _GEN_120 = io_rd_id == 12'h3b2 ? mhartid : _GEN_115; // @[regs.scala 286:42 regs.scala 68:30]
  wire [63:0] _GEN_121 = io_rd_id == 12'h3b1 ? _pmpaddr0_T : pmpaddr1; // @[regs.scala 284:42 regs.scala 285:18 regs.scala 63:30]
  wire [63:0] _GEN_122 = io_rd_id == 12'h3b1 ? pmpaddr2 : _GEN_116; // @[regs.scala 284:42 regs.scala 64:30]
  wire [63:0] _GEN_123 = io_rd_id == 12'h3b1 ? pmpaddr3 : _GEN_117; // @[regs.scala 284:42 regs.scala 65:30]
  wire [63:0] _GEN_125 = io_rd_id == 12'h3b1 ? uscratch : _GEN_119; // @[regs.scala 284:42 regs.scala 66:30]
  wire [63:0] _GEN_126 = io_rd_id == 12'h3b1 ? mhartid : _GEN_120; // @[regs.scala 284:42 regs.scala 68:30]
  wire [63:0] _GEN_127 = io_rd_id == 12'h3b0 ? _pmpaddr0_T : pmpaddr0; // @[regs.scala 282:42 regs.scala 283:18 regs.scala 62:30]
  wire [63:0] _GEN_128 = io_rd_id == 12'h3b0 ? pmpaddr1 : _GEN_121; // @[regs.scala 282:42 regs.scala 63:30]
  wire [63:0] _GEN_129 = io_rd_id == 12'h3b0 ? pmpaddr2 : _GEN_122; // @[regs.scala 282:42 regs.scala 64:30]
  wire [63:0] _GEN_130 = io_rd_id == 12'h3b0 ? pmpaddr3 : _GEN_123; // @[regs.scala 282:42 regs.scala 65:30]
  wire [63:0] _GEN_132 = io_rd_id == 12'h3b0 ? uscratch : _GEN_125; // @[regs.scala 282:42 regs.scala 66:30]
  wire [63:0] _GEN_133 = io_rd_id == 12'h3b0 ? mhartid : _GEN_126; // @[regs.scala 282:42 regs.scala 68:30]
  wire [63:0] _GEN_134 = io_rd_id == 12'h144 ? _mip_T_36 : _GEN_47; // @[regs.scala 280:37 regs.scala 281:13]
  wire [63:0] _GEN_135 = io_rd_id == 12'h144 ? pmpaddr0 : _GEN_127; // @[regs.scala 280:37 regs.scala 62:30]
  wire [63:0] _GEN_136 = io_rd_id == 12'h144 ? pmpaddr1 : _GEN_128; // @[regs.scala 280:37 regs.scala 63:30]
  wire [63:0] _GEN_137 = io_rd_id == 12'h144 ? pmpaddr2 : _GEN_129; // @[regs.scala 280:37 regs.scala 64:30]
  wire [63:0] _GEN_138 = io_rd_id == 12'h144 ? pmpaddr3 : _GEN_130; // @[regs.scala 280:37 regs.scala 65:30]
  wire [63:0] _GEN_140 = io_rd_id == 12'h144 ? uscratch : _GEN_132; // @[regs.scala 280:37 regs.scala 66:30]
  wire [63:0] _GEN_141 = io_rd_id == 12'h144 ? mhartid : _GEN_133; // @[regs.scala 280:37 regs.scala 68:30]
  wire [63:0] _GEN_142 = io_rd_id == 12'h104 ? _mie_T_3 : mie; // @[regs.scala 278:37 regs.scala 279:13 regs.scala 50:30]
  wire [63:0] _GEN_143 = io_rd_id == 12'h104 ? _GEN_47 : _GEN_134; // @[regs.scala 278:37]
  wire [63:0] _GEN_144 = io_rd_id == 12'h104 ? pmpaddr0 : _GEN_135; // @[regs.scala 278:37 regs.scala 62:30]
  wire [63:0] _GEN_145 = io_rd_id == 12'h104 ? pmpaddr1 : _GEN_136; // @[regs.scala 278:37 regs.scala 63:30]
  wire [63:0] _GEN_146 = io_rd_id == 12'h104 ? pmpaddr2 : _GEN_137; // @[regs.scala 278:37 regs.scala 64:30]
  wire [63:0] _GEN_147 = io_rd_id == 12'h104 ? pmpaddr3 : _GEN_138; // @[regs.scala 278:37 regs.scala 65:30]
  wire [63:0] _GEN_149 = io_rd_id == 12'h104 ? uscratch : _GEN_140; // @[regs.scala 278:37 regs.scala 66:30]
  wire [63:0] _GEN_150 = io_rd_id == 12'h104 ? mhartid : _GEN_141; // @[regs.scala 278:37 regs.scala 68:30]
  wire [63:0] _GEN_151 = io_rd_id == 12'h100 ? _mstatus_T_14 : _GEN_33; // @[regs.scala 274:41 regs.scala 277:17]
  wire [63:0] _GEN_152 = io_rd_id == 12'h100 ? mie : _GEN_142; // @[regs.scala 274:41 regs.scala 50:30]
  wire [63:0] _GEN_153 = io_rd_id == 12'h100 ? _GEN_47 : _GEN_143; // @[regs.scala 274:41]
  wire [63:0] _GEN_154 = io_rd_id == 12'h100 ? pmpaddr0 : _GEN_144; // @[regs.scala 274:41 regs.scala 62:30]
  wire [63:0] _GEN_155 = io_rd_id == 12'h100 ? pmpaddr1 : _GEN_145; // @[regs.scala 274:41 regs.scala 63:30]
  wire [63:0] _GEN_156 = io_rd_id == 12'h100 ? pmpaddr2 : _GEN_146; // @[regs.scala 274:41 regs.scala 64:30]
  wire [63:0] _GEN_157 = io_rd_id == 12'h100 ? pmpaddr3 : _GEN_147; // @[regs.scala 274:41 regs.scala 65:30]
  wire [63:0] _GEN_159 = io_rd_id == 12'h100 ? uscratch : _GEN_149; // @[regs.scala 274:41 regs.scala 66:30]
  wire [63:0] _GEN_160 = io_rd_id == 12'h100 ? mhartid : _GEN_150; // @[regs.scala 274:41 regs.scala 68:30]
  wire [63:0] _GEN_161 = io_rd_id == 12'h142 ? io_rd_data : _GEN_34; // @[regs.scala 272:40 regs.scala 273:16]
  wire [63:0] _GEN_162 = io_rd_id == 12'h142 ? _GEN_33 : _GEN_151; // @[regs.scala 272:40]
  wire [63:0] _GEN_163 = io_rd_id == 12'h142 ? mie : _GEN_152; // @[regs.scala 272:40 regs.scala 50:30]
  wire [63:0] _GEN_164 = io_rd_id == 12'h142 ? _GEN_47 : _GEN_153; // @[regs.scala 272:40]
  wire [63:0] _GEN_165 = io_rd_id == 12'h142 ? pmpaddr0 : _GEN_154; // @[regs.scala 272:40 regs.scala 62:30]
  wire [63:0] _GEN_166 = io_rd_id == 12'h142 ? pmpaddr1 : _GEN_155; // @[regs.scala 272:40 regs.scala 63:30]
  wire [63:0] _GEN_167 = io_rd_id == 12'h142 ? pmpaddr2 : _GEN_156; // @[regs.scala 272:40 regs.scala 64:30]
  wire [63:0] _GEN_168 = io_rd_id == 12'h142 ? pmpaddr3 : _GEN_157; // @[regs.scala 272:40 regs.scala 65:30]
  wire [63:0] _GEN_170 = io_rd_id == 12'h142 ? uscratch : _GEN_159; // @[regs.scala 272:40 regs.scala 66:30]
  wire [63:0] _GEN_171 = io_rd_id == 12'h142 ? mhartid : _GEN_160; // @[regs.scala 272:40 regs.scala 68:30]
  wire [63:0] _GEN_172 = io_rd_id == 12'h180 ? _satp_T_3 : satp; // @[regs.scala 270:38 regs.scala 271:14 regs.scala 60:30]
  wire [63:0] _GEN_173 = io_rd_id == 12'h180 ? _GEN_34 : _GEN_161; // @[regs.scala 270:38]
  wire [63:0] _GEN_174 = io_rd_id == 12'h180 ? _GEN_33 : _GEN_162; // @[regs.scala 270:38]
  wire [63:0] _GEN_175 = io_rd_id == 12'h180 ? mie : _GEN_163; // @[regs.scala 270:38 regs.scala 50:30]
  wire [63:0] _GEN_176 = io_rd_id == 12'h180 ? _GEN_47 : _GEN_164; // @[regs.scala 270:38]
  wire [63:0] _GEN_177 = io_rd_id == 12'h180 ? pmpaddr0 : _GEN_165; // @[regs.scala 270:38 regs.scala 62:30]
  wire [63:0] _GEN_178 = io_rd_id == 12'h180 ? pmpaddr1 : _GEN_166; // @[regs.scala 270:38 regs.scala 63:30]
  wire [63:0] _GEN_179 = io_rd_id == 12'h180 ? pmpaddr2 : _GEN_167; // @[regs.scala 270:38 regs.scala 64:30]
  wire [63:0] _GEN_180 = io_rd_id == 12'h180 ? pmpaddr3 : _GEN_168; // @[regs.scala 270:38 regs.scala 65:30]
  wire [63:0] _GEN_182 = io_rd_id == 12'h180 ? uscratch : _GEN_170; // @[regs.scala 270:38 regs.scala 66:30]
  wire [63:0] _GEN_183 = io_rd_id == 12'h180 ? mhartid : _GEN_171; // @[regs.scala 270:38 regs.scala 68:30]
  wire [63:0] _GEN_184 = io_rd_id == 12'h105 ? io_rd_data : stvec; // @[regs.scala 268:39 regs.scala 269:15 regs.scala 59:30]
  wire [63:0] _GEN_185 = io_rd_id == 12'h105 ? satp : _GEN_172; // @[regs.scala 268:39 regs.scala 60:30]
  wire [63:0] _GEN_186 = io_rd_id == 12'h105 ? _GEN_34 : _GEN_173; // @[regs.scala 268:39]
  wire [63:0] _GEN_187 = io_rd_id == 12'h105 ? _GEN_33 : _GEN_174; // @[regs.scala 268:39]
  wire [63:0] _GEN_188 = io_rd_id == 12'h105 ? mie : _GEN_175; // @[regs.scala 268:39 regs.scala 50:30]
  wire [63:0] _GEN_189 = io_rd_id == 12'h105 ? _GEN_47 : _GEN_176; // @[regs.scala 268:39]
  wire [63:0] _GEN_190 = io_rd_id == 12'h105 ? pmpaddr0 : _GEN_177; // @[regs.scala 268:39 regs.scala 62:30]
  wire [63:0] _GEN_191 = io_rd_id == 12'h105 ? pmpaddr1 : _GEN_178; // @[regs.scala 268:39 regs.scala 63:30]
  wire [63:0] _GEN_192 = io_rd_id == 12'h105 ? pmpaddr2 : _GEN_179; // @[regs.scala 268:39 regs.scala 64:30]
  wire [63:0] _GEN_193 = io_rd_id == 12'h105 ? pmpaddr3 : _GEN_180; // @[regs.scala 268:39 regs.scala 65:30]
  wire [63:0] _GEN_195 = io_rd_id == 12'h105 ? uscratch : _GEN_182; // @[regs.scala 268:39 regs.scala 66:30]
  wire [63:0] _GEN_196 = io_rd_id == 12'h105 ? mhartid : _GEN_183; // @[regs.scala 268:39 regs.scala 68:30]
  wire [63:0] _GEN_197 = io_rd_id == 12'h140 ? io_rd_data : sscratch; // @[regs.scala 266:42 regs.scala 267:18 regs.scala 58:30]
  wire [63:0] _GEN_198 = io_rd_id == 12'h140 ? stvec : _GEN_184; // @[regs.scala 266:42 regs.scala 59:30]
  wire [63:0] _GEN_199 = io_rd_id == 12'h140 ? satp : _GEN_185; // @[regs.scala 266:42 regs.scala 60:30]
  wire [63:0] _GEN_200 = io_rd_id == 12'h140 ? _GEN_34 : _GEN_186; // @[regs.scala 266:42]
  wire [63:0] _GEN_201 = io_rd_id == 12'h140 ? _GEN_33 : _GEN_187; // @[regs.scala 266:42]
  wire [63:0] _GEN_202 = io_rd_id == 12'h140 ? mie : _GEN_188; // @[regs.scala 266:42 regs.scala 50:30]
  wire [63:0] _GEN_203 = io_rd_id == 12'h140 ? _GEN_47 : _GEN_189; // @[regs.scala 266:42]
  wire [63:0] _GEN_204 = io_rd_id == 12'h140 ? pmpaddr0 : _GEN_190; // @[regs.scala 266:42 regs.scala 62:30]
  wire [63:0] _GEN_205 = io_rd_id == 12'h140 ? pmpaddr1 : _GEN_191; // @[regs.scala 266:42 regs.scala 63:30]
  wire [63:0] _GEN_206 = io_rd_id == 12'h140 ? pmpaddr2 : _GEN_192; // @[regs.scala 266:42 regs.scala 64:30]
  wire [63:0] _GEN_207 = io_rd_id == 12'h140 ? pmpaddr3 : _GEN_193; // @[regs.scala 266:42 regs.scala 65:30]
  wire [63:0] _GEN_209 = io_rd_id == 12'h140 ? uscratch : _GEN_195; // @[regs.scala 266:42 regs.scala 66:30]
  wire [63:0] _GEN_210 = io_rd_id == 12'h140 ? mhartid : _GEN_196; // @[regs.scala 266:42 regs.scala 68:30]
  wire [63:0] _GEN_211 = io_rd_id == 12'h143 ? io_rd_data : _GEN_36; // @[regs.scala 264:39 regs.scala 265:15]
  wire [63:0] _GEN_212 = io_rd_id == 12'h143 ? sscratch : _GEN_197; // @[regs.scala 264:39 regs.scala 58:30]
  wire [63:0] _GEN_213 = io_rd_id == 12'h143 ? stvec : _GEN_198; // @[regs.scala 264:39 regs.scala 59:30]
  wire [63:0] _GEN_214 = io_rd_id == 12'h143 ? satp : _GEN_199; // @[regs.scala 264:39 regs.scala 60:30]
  wire [63:0] _GEN_215 = io_rd_id == 12'h143 ? _GEN_34 : _GEN_200; // @[regs.scala 264:39]
  wire [63:0] _GEN_216 = io_rd_id == 12'h143 ? _GEN_33 : _GEN_201; // @[regs.scala 264:39]
  wire [63:0] _GEN_217 = io_rd_id == 12'h143 ? mie : _GEN_202; // @[regs.scala 264:39 regs.scala 50:30]
  wire [63:0] _GEN_218 = io_rd_id == 12'h143 ? _GEN_47 : _GEN_203; // @[regs.scala 264:39]
  wire [63:0] _GEN_219 = io_rd_id == 12'h143 ? pmpaddr0 : _GEN_204; // @[regs.scala 264:39 regs.scala 62:30]
  wire [63:0] _GEN_220 = io_rd_id == 12'h143 ? pmpaddr1 : _GEN_205; // @[regs.scala 264:39 regs.scala 63:30]
  wire [63:0] _GEN_221 = io_rd_id == 12'h143 ? pmpaddr2 : _GEN_206; // @[regs.scala 264:39 regs.scala 64:30]
  wire [63:0] _GEN_222 = io_rd_id == 12'h143 ? pmpaddr3 : _GEN_207; // @[regs.scala 264:39 regs.scala 65:30]
  wire [63:0] _GEN_224 = io_rd_id == 12'h143 ? uscratch : _GEN_209; // @[regs.scala 264:39 regs.scala 66:30]
  wire [63:0] _GEN_225 = io_rd_id == 12'h143 ? mhartid : _GEN_210; // @[regs.scala 264:39 regs.scala 68:30]
  wire [63:0] _GEN_226 = io_rd_id == 12'h141 ? io_rd_data : _GEN_35; // @[regs.scala 262:38 regs.scala 263:14]
  wire [63:0] _GEN_227 = io_rd_id == 12'h141 ? _GEN_36 : _GEN_211; // @[regs.scala 262:38]
  wire [63:0] _GEN_228 = io_rd_id == 12'h141 ? sscratch : _GEN_212; // @[regs.scala 262:38 regs.scala 58:30]
  wire [63:0] _GEN_229 = io_rd_id == 12'h141 ? stvec : _GEN_213; // @[regs.scala 262:38 regs.scala 59:30]
  wire [63:0] _GEN_230 = io_rd_id == 12'h141 ? satp : _GEN_214; // @[regs.scala 262:38 regs.scala 60:30]
  wire [63:0] _GEN_231 = io_rd_id == 12'h141 ? _GEN_34 : _GEN_215; // @[regs.scala 262:38]
  wire [63:0] _GEN_232 = io_rd_id == 12'h141 ? _GEN_33 : _GEN_216; // @[regs.scala 262:38]
  wire [63:0] _GEN_233 = io_rd_id == 12'h141 ? mie : _GEN_217; // @[regs.scala 262:38 regs.scala 50:30]
  wire [63:0] _GEN_234 = io_rd_id == 12'h141 ? _GEN_47 : _GEN_218; // @[regs.scala 262:38]
  wire [63:0] _GEN_235 = io_rd_id == 12'h141 ? pmpaddr0 : _GEN_219; // @[regs.scala 262:38 regs.scala 62:30]
  wire [63:0] _GEN_236 = io_rd_id == 12'h141 ? pmpaddr1 : _GEN_220; // @[regs.scala 262:38 regs.scala 63:30]
  wire [63:0] _GEN_237 = io_rd_id == 12'h141 ? pmpaddr2 : _GEN_221; // @[regs.scala 262:38 regs.scala 64:30]
  wire [63:0] _GEN_238 = io_rd_id == 12'h141 ? pmpaddr3 : _GEN_222; // @[regs.scala 262:38 regs.scala 65:30]
  wire [63:0] _GEN_240 = io_rd_id == 12'h141 ? uscratch : _GEN_224; // @[regs.scala 262:38 regs.scala 66:30]
  wire [63:0] _GEN_241 = io_rd_id == 12'h141 ? mhartid : _GEN_225; // @[regs.scala 262:38 regs.scala 68:30]
  wire [63:0] _GEN_242 = io_rd_id == 12'h106 ? io_rd_data : {{32'd0}, scounteren}; // @[regs.scala 260:44 regs.scala 261:20 regs.scala 55:30]
  wire [63:0] _GEN_243 = io_rd_id == 12'h106 ? _GEN_35 : _GEN_226; // @[regs.scala 260:44]
  wire [63:0] _GEN_244 = io_rd_id == 12'h106 ? _GEN_36 : _GEN_227; // @[regs.scala 260:44]
  wire [63:0] _GEN_245 = io_rd_id == 12'h106 ? sscratch : _GEN_228; // @[regs.scala 260:44 regs.scala 58:30]
  wire [63:0] _GEN_246 = io_rd_id == 12'h106 ? stvec : _GEN_229; // @[regs.scala 260:44 regs.scala 59:30]
  wire [63:0] _GEN_247 = io_rd_id == 12'h106 ? satp : _GEN_230; // @[regs.scala 260:44 regs.scala 60:30]
  wire [63:0] _GEN_248 = io_rd_id == 12'h106 ? _GEN_34 : _GEN_231; // @[regs.scala 260:44]
  wire [63:0] _GEN_249 = io_rd_id == 12'h106 ? _GEN_33 : _GEN_232; // @[regs.scala 260:44]
  wire [63:0] _GEN_250 = io_rd_id == 12'h106 ? mie : _GEN_233; // @[regs.scala 260:44 regs.scala 50:30]
  wire [63:0] _GEN_251 = io_rd_id == 12'h106 ? _GEN_47 : _GEN_234; // @[regs.scala 260:44]
  wire [63:0] _GEN_252 = io_rd_id == 12'h106 ? pmpaddr0 : _GEN_235; // @[regs.scala 260:44 regs.scala 62:30]
  wire [63:0] _GEN_253 = io_rd_id == 12'h106 ? pmpaddr1 : _GEN_236; // @[regs.scala 260:44 regs.scala 63:30]
  wire [63:0] _GEN_254 = io_rd_id == 12'h106 ? pmpaddr2 : _GEN_237; // @[regs.scala 260:44 regs.scala 64:30]
  wire [63:0] _GEN_255 = io_rd_id == 12'h106 ? pmpaddr3 : _GEN_238; // @[regs.scala 260:44 regs.scala 65:30]
  wire [63:0] _GEN_257 = io_rd_id == 12'h106 ? uscratch : _GEN_240; // @[regs.scala 260:44 regs.scala 66:30]
  wire [63:0] _GEN_258 = io_rd_id == 12'h106 ? mhartid : _GEN_241; // @[regs.scala 260:44 regs.scala 68:30]
  wire [63:0] _GEN_259 = io_rd_id == 12'h306 ? io_rd_data : {{32'd0}, mcounteren}; // @[regs.scala 258:44 regs.scala 259:20 regs.scala 54:30]
  wire [63:0] _GEN_260 = io_rd_id == 12'h306 ? {{32'd0}, scounteren} : _GEN_242; // @[regs.scala 258:44 regs.scala 55:30]
  wire [63:0] _GEN_261 = io_rd_id == 12'h306 ? _GEN_35 : _GEN_243; // @[regs.scala 258:44]
  wire [63:0] _GEN_262 = io_rd_id == 12'h306 ? _GEN_36 : _GEN_244; // @[regs.scala 258:44]
  wire [63:0] _GEN_263 = io_rd_id == 12'h306 ? sscratch : _GEN_245; // @[regs.scala 258:44 regs.scala 58:30]
  wire [63:0] _GEN_264 = io_rd_id == 12'h306 ? stvec : _GEN_246; // @[regs.scala 258:44 regs.scala 59:30]
  wire [63:0] _GEN_265 = io_rd_id == 12'h306 ? satp : _GEN_247; // @[regs.scala 258:44 regs.scala 60:30]
  wire [63:0] _GEN_266 = io_rd_id == 12'h306 ? _GEN_34 : _GEN_248; // @[regs.scala 258:44]
  wire [63:0] _GEN_267 = io_rd_id == 12'h306 ? _GEN_33 : _GEN_249; // @[regs.scala 258:44]
  wire [63:0] _GEN_268 = io_rd_id == 12'h306 ? mie : _GEN_250; // @[regs.scala 258:44 regs.scala 50:30]
  wire [63:0] _GEN_269 = io_rd_id == 12'h306 ? _GEN_47 : _GEN_251; // @[regs.scala 258:44]
  wire [63:0] _GEN_270 = io_rd_id == 12'h306 ? pmpaddr0 : _GEN_252; // @[regs.scala 258:44 regs.scala 62:30]
  wire [63:0] _GEN_271 = io_rd_id == 12'h306 ? pmpaddr1 : _GEN_253; // @[regs.scala 258:44 regs.scala 63:30]
  wire [63:0] _GEN_272 = io_rd_id == 12'h306 ? pmpaddr2 : _GEN_254; // @[regs.scala 258:44 regs.scala 64:30]
  wire [63:0] _GEN_273 = io_rd_id == 12'h306 ? pmpaddr3 : _GEN_255; // @[regs.scala 258:44 regs.scala 65:30]
  wire [63:0] _GEN_275 = io_rd_id == 12'h306 ? uscratch : _GEN_257; // @[regs.scala 258:44 regs.scala 66:30]
  wire [63:0] _GEN_276 = io_rd_id == 12'h306 ? mhartid : _GEN_258; // @[regs.scala 258:44 regs.scala 68:30]
  wire [63:0] _GEN_277 = io_rd_id == 12'h303 ? _mideleg_T : mideleg; // @[regs.scala 256:41 regs.scala 257:17 regs.scala 53:30]
  wire [63:0] _GEN_278 = io_rd_id == 12'h303 ? {{32'd0}, mcounteren} : _GEN_259; // @[regs.scala 256:41 regs.scala 54:30]
  wire [63:0] _GEN_279 = io_rd_id == 12'h303 ? {{32'd0}, scounteren} : _GEN_260; // @[regs.scala 256:41 regs.scala 55:30]
  wire [63:0] _GEN_280 = io_rd_id == 12'h303 ? _GEN_35 : _GEN_261; // @[regs.scala 256:41]
  wire [63:0] _GEN_281 = io_rd_id == 12'h303 ? _GEN_36 : _GEN_262; // @[regs.scala 256:41]
  wire [63:0] _GEN_282 = io_rd_id == 12'h303 ? sscratch : _GEN_263; // @[regs.scala 256:41 regs.scala 58:30]
  wire [63:0] _GEN_283 = io_rd_id == 12'h303 ? stvec : _GEN_264; // @[regs.scala 256:41 regs.scala 59:30]
  wire [63:0] _GEN_284 = io_rd_id == 12'h303 ? satp : _GEN_265; // @[regs.scala 256:41 regs.scala 60:30]
  wire [63:0] _GEN_285 = io_rd_id == 12'h303 ? _GEN_34 : _GEN_266; // @[regs.scala 256:41]
  wire [63:0] _GEN_286 = io_rd_id == 12'h303 ? _GEN_33 : _GEN_267; // @[regs.scala 256:41]
  wire [63:0] _GEN_287 = io_rd_id == 12'h303 ? mie : _GEN_268; // @[regs.scala 256:41 regs.scala 50:30]
  wire [63:0] _GEN_288 = io_rd_id == 12'h303 ? _GEN_47 : _GEN_269; // @[regs.scala 256:41]
  wire [63:0] _GEN_289 = io_rd_id == 12'h303 ? pmpaddr0 : _GEN_270; // @[regs.scala 256:41 regs.scala 62:30]
  wire [63:0] _GEN_290 = io_rd_id == 12'h303 ? pmpaddr1 : _GEN_271; // @[regs.scala 256:41 regs.scala 63:30]
  wire [63:0] _GEN_291 = io_rd_id == 12'h303 ? pmpaddr2 : _GEN_272; // @[regs.scala 256:41 regs.scala 64:30]
  wire [63:0] _GEN_292 = io_rd_id == 12'h303 ? pmpaddr3 : _GEN_273; // @[regs.scala 256:41 regs.scala 65:30]
  wire [63:0] _GEN_294 = io_rd_id == 12'h303 ? uscratch : _GEN_275; // @[regs.scala 256:41 regs.scala 66:30]
  wire [63:0] _GEN_295 = io_rd_id == 12'h303 ? mhartid : _GEN_276; // @[regs.scala 256:41 regs.scala 68:30]
  wire [63:0] _GEN_296 = io_rd_id == 12'h302 ? _medeleg_T : medeleg; // @[regs.scala 254:41 regs.scala 255:17 regs.scala 52:30]
  wire [63:0] _GEN_297 = io_rd_id == 12'h302 ? mideleg : _GEN_277; // @[regs.scala 254:41 regs.scala 53:30]
  wire [63:0] _GEN_298 = io_rd_id == 12'h302 ? {{32'd0}, mcounteren} : _GEN_278; // @[regs.scala 254:41 regs.scala 54:30]
  wire [63:0] _GEN_299 = io_rd_id == 12'h302 ? {{32'd0}, scounteren} : _GEN_279; // @[regs.scala 254:41 regs.scala 55:30]
  wire [63:0] _GEN_300 = io_rd_id == 12'h302 ? _GEN_35 : _GEN_280; // @[regs.scala 254:41]
  wire [63:0] _GEN_301 = io_rd_id == 12'h302 ? _GEN_36 : _GEN_281; // @[regs.scala 254:41]
  wire [63:0] _GEN_302 = io_rd_id == 12'h302 ? sscratch : _GEN_282; // @[regs.scala 254:41 regs.scala 58:30]
  wire [63:0] _GEN_303 = io_rd_id == 12'h302 ? stvec : _GEN_283; // @[regs.scala 254:41 regs.scala 59:30]
  wire [63:0] _GEN_304 = io_rd_id == 12'h302 ? satp : _GEN_284; // @[regs.scala 254:41 regs.scala 60:30]
  wire [63:0] _GEN_305 = io_rd_id == 12'h302 ? _GEN_34 : _GEN_285; // @[regs.scala 254:41]
  wire [63:0] _GEN_306 = io_rd_id == 12'h302 ? _GEN_33 : _GEN_286; // @[regs.scala 254:41]
  wire [63:0] _GEN_307 = io_rd_id == 12'h302 ? mie : _GEN_287; // @[regs.scala 254:41 regs.scala 50:30]
  wire [63:0] _GEN_308 = io_rd_id == 12'h302 ? _GEN_47 : _GEN_288; // @[regs.scala 254:41]
  wire [63:0] _GEN_309 = io_rd_id == 12'h302 ? pmpaddr0 : _GEN_289; // @[regs.scala 254:41 regs.scala 62:30]
  wire [63:0] _GEN_310 = io_rd_id == 12'h302 ? pmpaddr1 : _GEN_290; // @[regs.scala 254:41 regs.scala 63:30]
  wire [63:0] _GEN_311 = io_rd_id == 12'h302 ? pmpaddr2 : _GEN_291; // @[regs.scala 254:41 regs.scala 64:30]
  wire [63:0] _GEN_312 = io_rd_id == 12'h302 ? pmpaddr3 : _GEN_292; // @[regs.scala 254:41 regs.scala 65:30]
  wire [63:0] _GEN_314 = io_rd_id == 12'h302 ? uscratch : _GEN_294; // @[regs.scala 254:41 regs.scala 66:30]
  wire [63:0] _GEN_315 = io_rd_id == 12'h302 ? mhartid : _GEN_295; // @[regs.scala 254:41 regs.scala 68:30]
  wire [63:0] _GEN_316 = io_rd_id == 12'h342 ? io_rd_data : _GEN_37; // @[regs.scala 252:40 regs.scala 253:16]
  wire [63:0] _GEN_317 = io_rd_id == 12'h342 ? medeleg : _GEN_296; // @[regs.scala 252:40 regs.scala 52:30]
  wire [63:0] _GEN_318 = io_rd_id == 12'h342 ? mideleg : _GEN_297; // @[regs.scala 252:40 regs.scala 53:30]
  wire [63:0] _GEN_319 = io_rd_id == 12'h342 ? {{32'd0}, mcounteren} : _GEN_298; // @[regs.scala 252:40 regs.scala 54:30]
  wire [63:0] _GEN_320 = io_rd_id == 12'h342 ? {{32'd0}, scounteren} : _GEN_299; // @[regs.scala 252:40 regs.scala 55:30]
  wire [63:0] _GEN_321 = io_rd_id == 12'h342 ? _GEN_35 : _GEN_300; // @[regs.scala 252:40]
  wire [63:0] _GEN_322 = io_rd_id == 12'h342 ? _GEN_36 : _GEN_301; // @[regs.scala 252:40]
  wire [63:0] _GEN_323 = io_rd_id == 12'h342 ? sscratch : _GEN_302; // @[regs.scala 252:40 regs.scala 58:30]
  wire [63:0] _GEN_324 = io_rd_id == 12'h342 ? stvec : _GEN_303; // @[regs.scala 252:40 regs.scala 59:30]
  wire [63:0] _GEN_325 = io_rd_id == 12'h342 ? satp : _GEN_304; // @[regs.scala 252:40 regs.scala 60:30]
  wire [63:0] _GEN_326 = io_rd_id == 12'h342 ? _GEN_34 : _GEN_305; // @[regs.scala 252:40]
  wire [63:0] _GEN_327 = io_rd_id == 12'h342 ? _GEN_33 : _GEN_306; // @[regs.scala 252:40]
  wire [63:0] _GEN_328 = io_rd_id == 12'h342 ? mie : _GEN_307; // @[regs.scala 252:40 regs.scala 50:30]
  wire [63:0] _GEN_329 = io_rd_id == 12'h342 ? _GEN_47 : _GEN_308; // @[regs.scala 252:40]
  wire [63:0] _GEN_330 = io_rd_id == 12'h342 ? pmpaddr0 : _GEN_309; // @[regs.scala 252:40 regs.scala 62:30]
  wire [63:0] _GEN_331 = io_rd_id == 12'h342 ? pmpaddr1 : _GEN_310; // @[regs.scala 252:40 regs.scala 63:30]
  wire [63:0] _GEN_332 = io_rd_id == 12'h342 ? pmpaddr2 : _GEN_311; // @[regs.scala 252:40 regs.scala 64:30]
  wire [63:0] _GEN_333 = io_rd_id == 12'h342 ? pmpaddr3 : _GEN_312; // @[regs.scala 252:40 regs.scala 65:30]
  wire [63:0] _GEN_335 = io_rd_id == 12'h342 ? uscratch : _GEN_314; // @[regs.scala 252:40 regs.scala 66:30]
  wire [63:0] _GEN_336 = io_rd_id == 12'h342 ? mhartid : _GEN_315; // @[regs.scala 252:40 regs.scala 68:30]
  wire [63:0] _GEN_337 = io_rd_id == 12'h344 ? _mip_T_32 : _GEN_329; // @[regs.scala 250:37 regs.scala 251:13]
  wire [63:0] _GEN_338 = io_rd_id == 12'h344 ? _GEN_37 : _GEN_316; // @[regs.scala 250:37]
  wire [63:0] _GEN_339 = io_rd_id == 12'h344 ? medeleg : _GEN_317; // @[regs.scala 250:37 regs.scala 52:30]
  wire [63:0] _GEN_340 = io_rd_id == 12'h344 ? mideleg : _GEN_318; // @[regs.scala 250:37 regs.scala 53:30]
  wire [63:0] _GEN_341 = io_rd_id == 12'h344 ? {{32'd0}, mcounteren} : _GEN_319; // @[regs.scala 250:37 regs.scala 54:30]
  wire [63:0] _GEN_342 = io_rd_id == 12'h344 ? {{32'd0}, scounteren} : _GEN_320; // @[regs.scala 250:37 regs.scala 55:30]
  wire [63:0] _GEN_343 = io_rd_id == 12'h344 ? _GEN_35 : _GEN_321; // @[regs.scala 250:37]
  wire [63:0] _GEN_344 = io_rd_id == 12'h344 ? _GEN_36 : _GEN_322; // @[regs.scala 250:37]
  wire [63:0] _GEN_345 = io_rd_id == 12'h344 ? sscratch : _GEN_323; // @[regs.scala 250:37 regs.scala 58:30]
  wire [63:0] _GEN_346 = io_rd_id == 12'h344 ? stvec : _GEN_324; // @[regs.scala 250:37 regs.scala 59:30]
  wire [63:0] _GEN_347 = io_rd_id == 12'h344 ? satp : _GEN_325; // @[regs.scala 250:37 regs.scala 60:30]
  wire [63:0] _GEN_348 = io_rd_id == 12'h344 ? _GEN_34 : _GEN_326; // @[regs.scala 250:37]
  wire [63:0] _GEN_349 = io_rd_id == 12'h344 ? _GEN_33 : _GEN_327; // @[regs.scala 250:37]
  wire [63:0] _GEN_350 = io_rd_id == 12'h344 ? mie : _GEN_328; // @[regs.scala 250:37 regs.scala 50:30]
  wire [63:0] _GEN_351 = io_rd_id == 12'h344 ? pmpaddr0 : _GEN_330; // @[regs.scala 250:37 regs.scala 62:30]
  wire [63:0] _GEN_352 = io_rd_id == 12'h344 ? pmpaddr1 : _GEN_331; // @[regs.scala 250:37 regs.scala 63:30]
  wire [63:0] _GEN_353 = io_rd_id == 12'h344 ? pmpaddr2 : _GEN_332; // @[regs.scala 250:37 regs.scala 64:30]
  wire [63:0] _GEN_354 = io_rd_id == 12'h344 ? pmpaddr3 : _GEN_333; // @[regs.scala 250:37 regs.scala 65:30]
  wire [63:0] _GEN_356 = io_rd_id == 12'h344 ? uscratch : _GEN_335; // @[regs.scala 250:37 regs.scala 66:30]
  wire [63:0] _GEN_357 = io_rd_id == 12'h344 ? mhartid : _GEN_336; // @[regs.scala 250:37 regs.scala 68:30]
  wire [63:0] _GEN_358 = io_rd_id == 12'h304 ? io_rd_data : _GEN_350; // @[regs.scala 248:37 regs.scala 249:13]
  wire [63:0] _GEN_359 = io_rd_id == 12'h304 ? _GEN_47 : _GEN_337; // @[regs.scala 248:37]
  wire [63:0] _GEN_360 = io_rd_id == 12'h304 ? _GEN_37 : _GEN_338; // @[regs.scala 248:37]
  wire [63:0] _GEN_361 = io_rd_id == 12'h304 ? medeleg : _GEN_339; // @[regs.scala 248:37 regs.scala 52:30]
  wire [63:0] _GEN_362 = io_rd_id == 12'h304 ? mideleg : _GEN_340; // @[regs.scala 248:37 regs.scala 53:30]
  wire [63:0] _GEN_363 = io_rd_id == 12'h304 ? {{32'd0}, mcounteren} : _GEN_341; // @[regs.scala 248:37 regs.scala 54:30]
  wire [63:0] _GEN_364 = io_rd_id == 12'h304 ? {{32'd0}, scounteren} : _GEN_342; // @[regs.scala 248:37 regs.scala 55:30]
  wire [63:0] _GEN_365 = io_rd_id == 12'h304 ? _GEN_35 : _GEN_343; // @[regs.scala 248:37]
  wire [63:0] _GEN_366 = io_rd_id == 12'h304 ? _GEN_36 : _GEN_344; // @[regs.scala 248:37]
  wire [63:0] _GEN_367 = io_rd_id == 12'h304 ? sscratch : _GEN_345; // @[regs.scala 248:37 regs.scala 58:30]
  wire [63:0] _GEN_368 = io_rd_id == 12'h304 ? stvec : _GEN_346; // @[regs.scala 248:37 regs.scala 59:30]
  wire [63:0] _GEN_369 = io_rd_id == 12'h304 ? satp : _GEN_347; // @[regs.scala 248:37 regs.scala 60:30]
  wire [63:0] _GEN_370 = io_rd_id == 12'h304 ? _GEN_34 : _GEN_348; // @[regs.scala 248:37]
  wire [63:0] _GEN_371 = io_rd_id == 12'h304 ? _GEN_33 : _GEN_349; // @[regs.scala 248:37]
  wire [63:0] _GEN_372 = io_rd_id == 12'h304 ? pmpaddr0 : _GEN_351; // @[regs.scala 248:37 regs.scala 62:30]
  wire [63:0] _GEN_373 = io_rd_id == 12'h304 ? pmpaddr1 : _GEN_352; // @[regs.scala 248:37 regs.scala 63:30]
  wire [63:0] _GEN_374 = io_rd_id == 12'h304 ? pmpaddr2 : _GEN_353; // @[regs.scala 248:37 regs.scala 64:30]
  wire [63:0] _GEN_375 = io_rd_id == 12'h304 ? pmpaddr3 : _GEN_354; // @[regs.scala 248:37 regs.scala 65:30]
  wire [63:0] _GEN_377 = io_rd_id == 12'h304 ? uscratch : _GEN_356; // @[regs.scala 248:37 regs.scala 66:30]
  wire [63:0] _GEN_378 = io_rd_id == 12'h304 ? mhartid : _GEN_357; // @[regs.scala 248:37 regs.scala 68:30]
  wire [63:0] _GEN_379 = io_rd_id == 12'h305 ? io_rd_data : mtvec; // @[regs.scala 246:39 regs.scala 247:15 regs.scala 49:30]
  wire [63:0] _GEN_380 = io_rd_id == 12'h305 ? mie : _GEN_358; // @[regs.scala 246:39 regs.scala 50:30]
  wire [63:0] _GEN_381 = io_rd_id == 12'h305 ? _GEN_47 : _GEN_359; // @[regs.scala 246:39]
  wire [63:0] _GEN_382 = io_rd_id == 12'h305 ? _GEN_37 : _GEN_360; // @[regs.scala 246:39]
  wire [63:0] _GEN_383 = io_rd_id == 12'h305 ? medeleg : _GEN_361; // @[regs.scala 246:39 regs.scala 52:30]
  wire [63:0] _GEN_384 = io_rd_id == 12'h305 ? mideleg : _GEN_362; // @[regs.scala 246:39 regs.scala 53:30]
  wire [63:0] _GEN_385 = io_rd_id == 12'h305 ? {{32'd0}, mcounteren} : _GEN_363; // @[regs.scala 246:39 regs.scala 54:30]
  wire [63:0] _GEN_386 = io_rd_id == 12'h305 ? {{32'd0}, scounteren} : _GEN_364; // @[regs.scala 246:39 regs.scala 55:30]
  wire [63:0] _GEN_387 = io_rd_id == 12'h305 ? _GEN_35 : _GEN_365; // @[regs.scala 246:39]
  wire [63:0] _GEN_388 = io_rd_id == 12'h305 ? _GEN_36 : _GEN_366; // @[regs.scala 246:39]
  wire [63:0] _GEN_389 = io_rd_id == 12'h305 ? sscratch : _GEN_367; // @[regs.scala 246:39 regs.scala 58:30]
  wire [63:0] _GEN_390 = io_rd_id == 12'h305 ? stvec : _GEN_368; // @[regs.scala 246:39 regs.scala 59:30]
  wire [63:0] _GEN_391 = io_rd_id == 12'h305 ? satp : _GEN_369; // @[regs.scala 246:39 regs.scala 60:30]
  wire [63:0] _GEN_392 = io_rd_id == 12'h305 ? _GEN_34 : _GEN_370; // @[regs.scala 246:39]
  wire [63:0] _GEN_393 = io_rd_id == 12'h305 ? _GEN_33 : _GEN_371; // @[regs.scala 246:39]
  wire [63:0] _GEN_394 = io_rd_id == 12'h305 ? pmpaddr0 : _GEN_372; // @[regs.scala 246:39 regs.scala 62:30]
  wire [63:0] _GEN_395 = io_rd_id == 12'h305 ? pmpaddr1 : _GEN_373; // @[regs.scala 246:39 regs.scala 63:30]
  wire [63:0] _GEN_396 = io_rd_id == 12'h305 ? pmpaddr2 : _GEN_374; // @[regs.scala 246:39 regs.scala 64:30]
  wire [63:0] _GEN_397 = io_rd_id == 12'h305 ? pmpaddr3 : _GEN_375; // @[regs.scala 246:39 regs.scala 65:30]
  wire [63:0] _GEN_399 = io_rd_id == 12'h305 ? uscratch : _GEN_377; // @[regs.scala 246:39 regs.scala 66:30]
  wire [63:0] _GEN_400 = io_rd_id == 12'h305 ? mhartid : _GEN_378; // @[regs.scala 246:39 regs.scala 68:30]
  wire [63:0] _GEN_401 = io_rd_id == 12'h340 ? io_rd_data : mscratch; // @[regs.scala 244:42 regs.scala 245:18 regs.scala 47:30]
  wire [63:0] _GEN_402 = io_rd_id == 12'h340 ? mtvec : _GEN_379; // @[regs.scala 244:42 regs.scala 49:30]
  wire [63:0] _GEN_403 = io_rd_id == 12'h340 ? mie : _GEN_380; // @[regs.scala 244:42 regs.scala 50:30]
  wire [63:0] _GEN_404 = io_rd_id == 12'h340 ? _GEN_47 : _GEN_381; // @[regs.scala 244:42]
  wire [63:0] _GEN_405 = io_rd_id == 12'h340 ? _GEN_37 : _GEN_382; // @[regs.scala 244:42]
  wire [63:0] _GEN_406 = io_rd_id == 12'h340 ? medeleg : _GEN_383; // @[regs.scala 244:42 regs.scala 52:30]
  wire [63:0] _GEN_407 = io_rd_id == 12'h340 ? mideleg : _GEN_384; // @[regs.scala 244:42 regs.scala 53:30]
  wire [63:0] _GEN_408 = io_rd_id == 12'h340 ? {{32'd0}, mcounteren} : _GEN_385; // @[regs.scala 244:42 regs.scala 54:30]
  wire [63:0] _GEN_409 = io_rd_id == 12'h340 ? {{32'd0}, scounteren} : _GEN_386; // @[regs.scala 244:42 regs.scala 55:30]
  wire [63:0] _GEN_410 = io_rd_id == 12'h340 ? _GEN_35 : _GEN_387; // @[regs.scala 244:42]
  wire [63:0] _GEN_411 = io_rd_id == 12'h340 ? _GEN_36 : _GEN_388; // @[regs.scala 244:42]
  wire [63:0] _GEN_412 = io_rd_id == 12'h340 ? sscratch : _GEN_389; // @[regs.scala 244:42 regs.scala 58:30]
  wire [63:0] _GEN_413 = io_rd_id == 12'h340 ? stvec : _GEN_390; // @[regs.scala 244:42 regs.scala 59:30]
  wire [63:0] _GEN_414 = io_rd_id == 12'h340 ? satp : _GEN_391; // @[regs.scala 244:42 regs.scala 60:30]
  wire [63:0] _GEN_415 = io_rd_id == 12'h340 ? _GEN_34 : _GEN_392; // @[regs.scala 244:42]
  wire [63:0] _GEN_416 = io_rd_id == 12'h340 ? _GEN_33 : _GEN_393; // @[regs.scala 244:42]
  wire [63:0] _GEN_417 = io_rd_id == 12'h340 ? pmpaddr0 : _GEN_394; // @[regs.scala 244:42 regs.scala 62:30]
  wire [63:0] _GEN_418 = io_rd_id == 12'h340 ? pmpaddr1 : _GEN_395; // @[regs.scala 244:42 regs.scala 63:30]
  wire [63:0] _GEN_419 = io_rd_id == 12'h340 ? pmpaddr2 : _GEN_396; // @[regs.scala 244:42 regs.scala 64:30]
  wire [63:0] _GEN_420 = io_rd_id == 12'h340 ? pmpaddr3 : _GEN_397; // @[regs.scala 244:42 regs.scala 65:30]
  wire [63:0] _GEN_422 = io_rd_id == 12'h340 ? uscratch : _GEN_399; // @[regs.scala 244:42 regs.scala 66:30]
  wire [63:0] _GEN_423 = io_rd_id == 12'h340 ? mhartid : _GEN_400; // @[regs.scala 244:42 regs.scala 68:30]
  wire [63:0] _GEN_424 = io_rd_id == 12'h343 ? io_rd_data : _GEN_39; // @[regs.scala 242:39 regs.scala 243:15]
  wire [63:0] _GEN_425 = io_rd_id == 12'h343 ? mscratch : _GEN_401; // @[regs.scala 242:39 regs.scala 47:30]
  wire [63:0] _GEN_426 = io_rd_id == 12'h343 ? mtvec : _GEN_402; // @[regs.scala 242:39 regs.scala 49:30]
  wire [63:0] _GEN_427 = io_rd_id == 12'h343 ? mie : _GEN_403; // @[regs.scala 242:39 regs.scala 50:30]
  wire [63:0] _GEN_428 = io_rd_id == 12'h343 ? _GEN_47 : _GEN_404; // @[regs.scala 242:39]
  wire [63:0] _GEN_429 = io_rd_id == 12'h343 ? _GEN_37 : _GEN_405; // @[regs.scala 242:39]
  wire [63:0] _GEN_430 = io_rd_id == 12'h343 ? medeleg : _GEN_406; // @[regs.scala 242:39 regs.scala 52:30]
  wire [63:0] _GEN_431 = io_rd_id == 12'h343 ? mideleg : _GEN_407; // @[regs.scala 242:39 regs.scala 53:30]
  wire [63:0] _GEN_432 = io_rd_id == 12'h343 ? {{32'd0}, mcounteren} : _GEN_408; // @[regs.scala 242:39 regs.scala 54:30]
  wire [63:0] _GEN_433 = io_rd_id == 12'h343 ? {{32'd0}, scounteren} : _GEN_409; // @[regs.scala 242:39 regs.scala 55:30]
  wire [63:0] _GEN_434 = io_rd_id == 12'h343 ? _GEN_35 : _GEN_410; // @[regs.scala 242:39]
  wire [63:0] _GEN_435 = io_rd_id == 12'h343 ? _GEN_36 : _GEN_411; // @[regs.scala 242:39]
  wire [63:0] _GEN_436 = io_rd_id == 12'h343 ? sscratch : _GEN_412; // @[regs.scala 242:39 regs.scala 58:30]
  wire [63:0] _GEN_437 = io_rd_id == 12'h343 ? stvec : _GEN_413; // @[regs.scala 242:39 regs.scala 59:30]
  wire [63:0] _GEN_438 = io_rd_id == 12'h343 ? satp : _GEN_414; // @[regs.scala 242:39 regs.scala 60:30]
  wire [63:0] _GEN_439 = io_rd_id == 12'h343 ? _GEN_34 : _GEN_415; // @[regs.scala 242:39]
  wire [63:0] _GEN_440 = io_rd_id == 12'h343 ? _GEN_33 : _GEN_416; // @[regs.scala 242:39]
  wire [63:0] _GEN_441 = io_rd_id == 12'h343 ? pmpaddr0 : _GEN_417; // @[regs.scala 242:39 regs.scala 62:30]
  wire [63:0] _GEN_442 = io_rd_id == 12'h343 ? pmpaddr1 : _GEN_418; // @[regs.scala 242:39 regs.scala 63:30]
  wire [63:0] _GEN_443 = io_rd_id == 12'h343 ? pmpaddr2 : _GEN_419; // @[regs.scala 242:39 regs.scala 64:30]
  wire [63:0] _GEN_444 = io_rd_id == 12'h343 ? pmpaddr3 : _GEN_420; // @[regs.scala 242:39 regs.scala 65:30]
  wire [63:0] _GEN_446 = io_rd_id == 12'h343 ? uscratch : _GEN_422; // @[regs.scala 242:39 regs.scala 66:30]
  wire [63:0] _GEN_447 = io_rd_id == 12'h343 ? mhartid : _GEN_423; // @[regs.scala 242:39 regs.scala 68:30]
  wire [63:0] _GEN_448 = io_rd_id == 12'h341 ? io_rd_data : _GEN_38; // @[regs.scala 240:38 regs.scala 241:14]
  wire [63:0] _GEN_449 = io_rd_id == 12'h341 ? _GEN_39 : _GEN_424; // @[regs.scala 240:38]
  wire [63:0] _GEN_450 = io_rd_id == 12'h341 ? mscratch : _GEN_425; // @[regs.scala 240:38 regs.scala 47:30]
  wire [63:0] _GEN_451 = io_rd_id == 12'h341 ? mtvec : _GEN_426; // @[regs.scala 240:38 regs.scala 49:30]
  wire [63:0] _GEN_452 = io_rd_id == 12'h341 ? mie : _GEN_427; // @[regs.scala 240:38 regs.scala 50:30]
  wire [63:0] _GEN_453 = io_rd_id == 12'h341 ? _GEN_47 : _GEN_428; // @[regs.scala 240:38]
  wire [63:0] _GEN_454 = io_rd_id == 12'h341 ? _GEN_37 : _GEN_429; // @[regs.scala 240:38]
  wire [63:0] _GEN_455 = io_rd_id == 12'h341 ? medeleg : _GEN_430; // @[regs.scala 240:38 regs.scala 52:30]
  wire [63:0] _GEN_456 = io_rd_id == 12'h341 ? mideleg : _GEN_431; // @[regs.scala 240:38 regs.scala 53:30]
  wire [63:0] _GEN_457 = io_rd_id == 12'h341 ? {{32'd0}, mcounteren} : _GEN_432; // @[regs.scala 240:38 regs.scala 54:30]
  wire [63:0] _GEN_458 = io_rd_id == 12'h341 ? {{32'd0}, scounteren} : _GEN_433; // @[regs.scala 240:38 regs.scala 55:30]
  wire [63:0] _GEN_459 = io_rd_id == 12'h341 ? _GEN_35 : _GEN_434; // @[regs.scala 240:38]
  wire [63:0] _GEN_460 = io_rd_id == 12'h341 ? _GEN_36 : _GEN_435; // @[regs.scala 240:38]
  wire [63:0] _GEN_461 = io_rd_id == 12'h341 ? sscratch : _GEN_436; // @[regs.scala 240:38 regs.scala 58:30]
  wire [63:0] _GEN_462 = io_rd_id == 12'h341 ? stvec : _GEN_437; // @[regs.scala 240:38 regs.scala 59:30]
  wire [63:0] _GEN_463 = io_rd_id == 12'h341 ? satp : _GEN_438; // @[regs.scala 240:38 regs.scala 60:30]
  wire [63:0] _GEN_464 = io_rd_id == 12'h341 ? _GEN_34 : _GEN_439; // @[regs.scala 240:38]
  wire [63:0] _GEN_465 = io_rd_id == 12'h341 ? _GEN_33 : _GEN_440; // @[regs.scala 240:38]
  wire [63:0] _GEN_466 = io_rd_id == 12'h341 ? pmpaddr0 : _GEN_441; // @[regs.scala 240:38 regs.scala 62:30]
  wire [63:0] _GEN_467 = io_rd_id == 12'h341 ? pmpaddr1 : _GEN_442; // @[regs.scala 240:38 regs.scala 63:30]
  wire [63:0] _GEN_468 = io_rd_id == 12'h341 ? pmpaddr2 : _GEN_443; // @[regs.scala 240:38 regs.scala 64:30]
  wire [63:0] _GEN_469 = io_rd_id == 12'h341 ? pmpaddr3 : _GEN_444; // @[regs.scala 240:38 regs.scala 65:30]
  wire [63:0] _GEN_471 = io_rd_id == 12'h341 ? uscratch : _GEN_446; // @[regs.scala 240:38 regs.scala 66:30]
  wire [63:0] _GEN_472 = io_rd_id == 12'h341 ? mhartid : _GEN_447; // @[regs.scala 240:38 regs.scala 68:30]
  wire [63:0] _GEN_483 = io_rd_id == 12'h300 ? {{32'd0}, mcounteren} : _GEN_457; // @[regs.scala 236:41 regs.scala 54:30]
  wire [63:0] _GEN_484 = io_rd_id == 12'h300 ? {{32'd0}, scounteren} : _GEN_458; // @[regs.scala 236:41 regs.scala 55:30]
  wire [63:0] _GEN_509 = io_rd_id == 12'h301 ? {{32'd0}, mcounteren} : _GEN_483; // @[regs.scala 234:38 regs.scala 54:30]
  wire [63:0] _GEN_510 = io_rd_id == 12'h301 ? {{32'd0}, scounteren} : _GEN_484; // @[regs.scala 234:38 regs.scala 55:30]
  wire [63:0] _GEN_535 = ~io_rd_en ? {{32'd0}, mcounteren} : _GEN_509; // @[regs.scala 233:20 regs.scala 54:30]
  wire [63:0] _GEN_536 = ~io_rd_en ? {{32'd0}, scounteren} : _GEN_510; // @[regs.scala 233:20 regs.scala 55:30]
  assign io_rs_data = io_rs_id == 12'h301 ? misa : _GEN_102; // @[regs.scala 171:32 regs.scala 172:20]
  assign io_rs_is_err = io_rs_id == 12'h301 ? 1'h0 : _GEN_103; // @[regs.scala 171:32 regs.scala 170:21]
  assign io_mmuState_priv = priv; // @[regs.scala 71:25]
  assign io_mmuState_mstatus = mstatus; // @[regs.scala 72:25]
  assign io_mmuState_satp = satp; // @[regs.scala 73:25]
  assign io_idState_priv = priv; // @[regs.scala 74:24]
  assign io_reg2if_seq_pc = forceJmp_seq_pc; // @[regs.scala 76:25]
  assign io_reg2if_valid = forceJmp_valid; // @[regs.scala 76:25]
  assign io_intr_out_en = intr_out_r_en; // @[regs.scala 125:17]
  assign io_intr_out_cause = intr_out_r_cause; // @[regs.scala 125:17]
  assign io_updateNextPc_seq_pc = forceJmp_seq_pc; // @[regs.scala 79:25]
  assign io_updateNextPc_valid = forceJmp_valid; // @[regs.scala 79:25]
  always @(posedge clock) begin
    if (reset) begin // @[regs.scala 42:30]
      priv <= 2'h3; // @[regs.scala 42:30]
    end else if (io_excep_en) begin // @[regs.scala 80:22]
      if (io_excep_etype == 2'h2) begin // @[regs.scala 81:44]
        priv <= _priv_T; // @[regs.scala 85:29]
      end else if (io_excep_etype == 2'h3) begin // @[regs.scala 88:50]
        priv <= mstatus[12:11]; // @[regs.scala 92:29]
      end else begin
        priv <= _GEN_6;
      end
    end
    if (reset) begin // @[regs.scala 43:30]
      misa <= 64'h800000000014112d; // @[regs.scala 43:30]
    end else if (!(~io_rd_en)) begin // @[regs.scala 233:20]
      if (io_rd_id == 12'h301) begin // @[regs.scala 234:38]
        misa <= io_rd_data; // @[regs.scala 235:14]
      end
    end
    if (reset) begin // @[regs.scala 44:30]
      mstatus <= 64'ha00000000; // @[regs.scala 44:30]
    end else if (~io_rd_en) begin // @[regs.scala 233:20]
      mstatus <= _GEN_33;
    end else if (io_rd_id == 12'h301) begin // @[regs.scala 234:38]
      mstatus <= _GEN_33;
    end else if (io_rd_id == 12'h300) begin // @[regs.scala 236:41]
      mstatus <= _mstatus_T_13; // @[regs.scala 239:17]
    end else begin
      mstatus <= _GEN_465;
    end
    if (reset) begin // @[regs.scala 45:30]
      mepc <= 64'h0; // @[regs.scala 45:30]
    end else if (~io_rd_en) begin // @[regs.scala 233:20]
      mepc <= _GEN_38;
    end else if (io_rd_id == 12'h301) begin // @[regs.scala 234:38]
      mepc <= _GEN_38;
    end else if (io_rd_id == 12'h300) begin // @[regs.scala 236:41]
      mepc <= _GEN_38;
    end else begin
      mepc <= _GEN_448;
    end
    if (reset) begin // @[regs.scala 46:30]
      mtval <= 64'h0; // @[regs.scala 46:30]
    end else if (~io_rd_en) begin // @[regs.scala 233:20]
      mtval <= _GEN_39;
    end else if (io_rd_id == 12'h301) begin // @[regs.scala 234:38]
      mtval <= _GEN_39;
    end else if (io_rd_id == 12'h300) begin // @[regs.scala 236:41]
      mtval <= _GEN_39;
    end else begin
      mtval <= _GEN_449;
    end
    if (reset) begin // @[regs.scala 47:30]
      mscratch <= 64'h0; // @[regs.scala 47:30]
    end else if (!(~io_rd_en)) begin // @[regs.scala 233:20]
      if (!(io_rd_id == 12'h301)) begin // @[regs.scala 234:38]
        if (!(io_rd_id == 12'h300)) begin // @[regs.scala 236:41]
          mscratch <= _GEN_450;
        end
      end
    end
    if (reset) begin // @[regs.scala 48:30]
      mcause <= 64'h0; // @[regs.scala 48:30]
    end else if (~io_rd_en) begin // @[regs.scala 233:20]
      mcause <= _GEN_37;
    end else if (io_rd_id == 12'h301) begin // @[regs.scala 234:38]
      mcause <= _GEN_37;
    end else if (io_rd_id == 12'h300) begin // @[regs.scala 236:41]
      mcause <= _GEN_37;
    end else begin
      mcause <= _GEN_454;
    end
    if (reset) begin // @[regs.scala 49:30]
      mtvec <= 64'h0; // @[regs.scala 49:30]
    end else if (!(~io_rd_en)) begin // @[regs.scala 233:20]
      if (!(io_rd_id == 12'h301)) begin // @[regs.scala 234:38]
        if (!(io_rd_id == 12'h300)) begin // @[regs.scala 236:41]
          mtvec <= _GEN_451;
        end
      end
    end
    if (reset) begin // @[regs.scala 50:30]
      mie <= 64'h0; // @[regs.scala 50:30]
    end else if (!(~io_rd_en)) begin // @[regs.scala 233:20]
      if (!(io_rd_id == 12'h301)) begin // @[regs.scala 234:38]
        if (!(io_rd_id == 12'h300)) begin // @[regs.scala 236:41]
          mie <= _GEN_452;
        end
      end
    end
    if (reset) begin // @[regs.scala 51:30]
      mip <= 64'h0; // @[regs.scala 51:30]
    end else if (~io_rd_en) begin // @[regs.scala 233:20]
      mip <= _GEN_47;
    end else if (io_rd_id == 12'h301) begin // @[regs.scala 234:38]
      mip <= _GEN_47;
    end else if (io_rd_id == 12'h300) begin // @[regs.scala 236:41]
      mip <= _GEN_47;
    end else begin
      mip <= _GEN_453;
    end
    if (reset) begin // @[regs.scala 52:30]
      medeleg <= 64'h0; // @[regs.scala 52:30]
    end else if (!(~io_rd_en)) begin // @[regs.scala 233:20]
      if (!(io_rd_id == 12'h301)) begin // @[regs.scala 234:38]
        if (!(io_rd_id == 12'h300)) begin // @[regs.scala 236:41]
          medeleg <= _GEN_455;
        end
      end
    end
    if (reset) begin // @[regs.scala 53:30]
      mideleg <= 64'h0; // @[regs.scala 53:30]
    end else if (!(~io_rd_en)) begin // @[regs.scala 233:20]
      if (!(io_rd_id == 12'h301)) begin // @[regs.scala 234:38]
        if (!(io_rd_id == 12'h300)) begin // @[regs.scala 236:41]
          mideleg <= _GEN_456;
        end
      end
    end
    if (reset) begin // @[regs.scala 54:30]
      mcounteren <= 32'h0; // @[regs.scala 54:30]
    end else begin
      mcounteren <= _GEN_535[31:0];
    end
    if (reset) begin // @[regs.scala 55:30]
      scounteren <= 32'h0; // @[regs.scala 55:30]
    end else begin
      scounteren <= _GEN_536[31:0];
    end
    if (reset) begin // @[regs.scala 56:30]
      sepc <= 64'h0; // @[regs.scala 56:30]
    end else if (~io_rd_en) begin // @[regs.scala 233:20]
      sepc <= _GEN_35;
    end else if (io_rd_id == 12'h301) begin // @[regs.scala 234:38]
      sepc <= _GEN_35;
    end else if (io_rd_id == 12'h300) begin // @[regs.scala 236:41]
      sepc <= _GEN_35;
    end else begin
      sepc <= _GEN_459;
    end
    if (reset) begin // @[regs.scala 57:30]
      stval <= 64'h0; // @[regs.scala 57:30]
    end else if (~io_rd_en) begin // @[regs.scala 233:20]
      stval <= _GEN_36;
    end else if (io_rd_id == 12'h301) begin // @[regs.scala 234:38]
      stval <= _GEN_36;
    end else if (io_rd_id == 12'h300) begin // @[regs.scala 236:41]
      stval <= _GEN_36;
    end else begin
      stval <= _GEN_460;
    end
    if (reset) begin // @[regs.scala 58:30]
      sscratch <= 64'h0; // @[regs.scala 58:30]
    end else if (!(~io_rd_en)) begin // @[regs.scala 233:20]
      if (!(io_rd_id == 12'h301)) begin // @[regs.scala 234:38]
        if (!(io_rd_id == 12'h300)) begin // @[regs.scala 236:41]
          sscratch <= _GEN_461;
        end
      end
    end
    if (reset) begin // @[regs.scala 59:30]
      stvec <= 64'h0; // @[regs.scala 59:30]
    end else if (!(~io_rd_en)) begin // @[regs.scala 233:20]
      if (!(io_rd_id == 12'h301)) begin // @[regs.scala 234:38]
        if (!(io_rd_id == 12'h300)) begin // @[regs.scala 236:41]
          stvec <= _GEN_462;
        end
      end
    end
    if (reset) begin // @[regs.scala 60:30]
      satp <= 64'h0; // @[regs.scala 60:30]
    end else if (!(~io_rd_en)) begin // @[regs.scala 233:20]
      if (!(io_rd_id == 12'h301)) begin // @[regs.scala 234:38]
        if (!(io_rd_id == 12'h300)) begin // @[regs.scala 236:41]
          satp <= _GEN_463;
        end
      end
    end
    if (reset) begin // @[regs.scala 61:30]
      scause <= 64'h0; // @[regs.scala 61:30]
    end else if (~io_rd_en) begin // @[regs.scala 233:20]
      scause <= _GEN_34;
    end else if (io_rd_id == 12'h301) begin // @[regs.scala 234:38]
      scause <= _GEN_34;
    end else if (io_rd_id == 12'h300) begin // @[regs.scala 236:41]
      scause <= _GEN_34;
    end else begin
      scause <= _GEN_464;
    end
    if (reset) begin // @[regs.scala 62:30]
      pmpaddr0 <= 64'h0; // @[regs.scala 62:30]
    end else if (!(~io_rd_en)) begin // @[regs.scala 233:20]
      if (!(io_rd_id == 12'h301)) begin // @[regs.scala 234:38]
        if (!(io_rd_id == 12'h300)) begin // @[regs.scala 236:41]
          pmpaddr0 <= _GEN_466;
        end
      end
    end
    if (reset) begin // @[regs.scala 63:30]
      pmpaddr1 <= 64'h0; // @[regs.scala 63:30]
    end else if (!(~io_rd_en)) begin // @[regs.scala 233:20]
      if (!(io_rd_id == 12'h301)) begin // @[regs.scala 234:38]
        if (!(io_rd_id == 12'h300)) begin // @[regs.scala 236:41]
          pmpaddr1 <= _GEN_467;
        end
      end
    end
    if (reset) begin // @[regs.scala 64:30]
      pmpaddr2 <= 64'h0; // @[regs.scala 64:30]
    end else if (!(~io_rd_en)) begin // @[regs.scala 233:20]
      if (!(io_rd_id == 12'h301)) begin // @[regs.scala 234:38]
        if (!(io_rd_id == 12'h300)) begin // @[regs.scala 236:41]
          pmpaddr2 <= _GEN_468;
        end
      end
    end
    if (reset) begin // @[regs.scala 65:30]
      pmpaddr3 <= 64'h0; // @[regs.scala 65:30]
    end else if (!(~io_rd_en)) begin // @[regs.scala 233:20]
      if (!(io_rd_id == 12'h301)) begin // @[regs.scala 234:38]
        if (!(io_rd_id == 12'h300)) begin // @[regs.scala 236:41]
          pmpaddr3 <= _GEN_469;
        end
      end
    end
    if (reset) begin // @[regs.scala 66:30]
      uscratch <= 64'h0; // @[regs.scala 66:30]
    end else if (!(~io_rd_en)) begin // @[regs.scala 233:20]
      if (!(io_rd_id == 12'h301)) begin // @[regs.scala 234:38]
        if (!(io_rd_id == 12'h300)) begin // @[regs.scala 236:41]
          uscratch <= _GEN_471;
        end
      end
    end
    if (reset) begin // @[regs.scala 68:30]
      mhartid <= 64'h0; // @[regs.scala 68:30]
    end else if (!(~io_rd_en)) begin // @[regs.scala 233:20]
      if (!(io_rd_id == 12'h301)) begin // @[regs.scala 234:38]
        if (!(io_rd_id == 12'h300)) begin // @[regs.scala 236:41]
          mhartid <= _GEN_472;
        end
      end
    end
    if (reset) begin // @[regs.scala 75:34]
      forceJmp_seq_pc <= 64'h0; // @[regs.scala 75:34]
    end else begin
      forceJmp_seq_pc <= _GEN_30[63:0];
    end
    if (reset) begin // @[regs.scala 75:34]
      forceJmp_valid <= 1'h0; // @[regs.scala 75:34]
    end else begin
      forceJmp_valid <= io_excep_en;
    end
    if (reset) begin // @[regs.scala 124:29]
      intr_out_r_en <= 1'h0; // @[regs.scala 124:29]
    end else begin
      intr_out_r_en <= enable_int != 64'h0; // @[regs.scala 158:19]
    end
    if (reset) begin // @[regs.scala 124:29]
      intr_out_r_cause <= 64'h0; // @[regs.scala 124:29]
    end else begin
      intr_out_r_cause <= _intr_out_r_cause_T_13; // @[regs.scala 160:22]
    end
    if (reset) begin // @[regs.scala 126:28]
      intr_seip <= 1'h0; // @[regs.scala 126:28]
    end else if (io_plic_s_clear) begin // @[regs.scala 142:26]
      intr_seip <= 1'h0; // @[regs.scala 143:19]
    end else begin
      intr_seip <= _GEN_44;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  priv = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  misa = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mstatus = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mepc = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mtval = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mscratch = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mcause = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  mtvec = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  mie = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  mip = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  medeleg = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mideleg = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  mcounteren = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  scounteren = _RAND_13[31:0];
  _RAND_14 = {2{`RANDOM}};
  sepc = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  stval = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  sscratch = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  stvec = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  satp = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  scause = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  pmpaddr0 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  pmpaddr1 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  pmpaddr2 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  pmpaddr3 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  uscratch = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  mhartid = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  forceJmp_seq_pc = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  forceJmp_valid = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  intr_out_r_en = _RAND_28[0:0];
  _RAND_29 = {2{`RANDOM}};
  intr_out_r_cause = _RAND_29[63:0];
  _RAND_30 = {1{`RANDOM}};
  intr_seip = _RAND_30[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 47:50]
  reg  state_1; // @[PRNG.scala 47:50]
  reg  state_2; // @[PRNG.scala 47:50]
  wire  _T = state_2 ^ state_1; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 69:10]
  assign io_out_1 = state_1; // @[PRNG.scala 69:10]
  assign io_out_2 = state_2; // @[PRNG.scala 69:10]
  always @(posedge clock) begin
    state_0 <= reset | _T; // @[PRNG.scala 47:50 PRNG.scala 47:50]
    if (reset) begin // @[PRNG.scala 47:50]
      state_1 <= 1'h0; // @[PRNG.scala 47:50]
    end else begin
      state_1 <= state_0;
    end
    if (reset) begin // @[PRNG.scala 47:50]
      state_2 <= 1'h0; // @[PRNG.scala 47:50]
    end else begin
      state_2 <= state_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_InstCache(
  input          clock,
  input          reset,
  input          io_instAxi_ra_ready,
  output         io_instAxi_ra_valid,
  output [31:0]  io_instAxi_ra_bits_addr,
  input          io_instAxi_rd_valid,
  input  [63:0]  io_instAxi_rd_bits_data,
  input          io_instAxi_rd_bits_last,
  input  [31:0]  io_icRead_addr,
  output [63:0]  io_icRead_inst,
  input          io_icRead_arvalid,
  output         io_icRead_ready,
  output         io_icRead_rvalid,
  input          io_flush,
  output [5:0]   io_ic2sr0_addr,
  output         io_ic2sr0_cen,
  output         io_ic2sr0_wen,
  output [127:0] io_ic2sr0_wmask,
  output [127:0] io_ic2sr0_wdata,
  input  [127:0] io_ic2sr0_rdata,
  output [5:0]   io_ic2sr1_addr,
  output         io_ic2sr1_cen,
  output         io_ic2sr1_wen,
  output [127:0] io_ic2sr1_wmask,
  output [127:0] io_ic2sr1_wdata,
  input  [127:0] io_ic2sr1_rdata,
  output [5:0]   io_ic2sr2_addr,
  output         io_ic2sr2_cen,
  output         io_ic2sr2_wen,
  output [127:0] io_ic2sr2_wmask,
  output [127:0] io_ic2sr2_wdata,
  input  [127:0] io_ic2sr2_rdata,
  output [5:0]   io_ic2sr3_addr,
  output         io_ic2sr3_cen,
  output         io_ic2sr3_wen,
  output [127:0] io_ic2sr3_wmask,
  output [127:0] io_ic2sr3_wdata,
  input  [127:0] io_ic2sr3_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
`endif // RANDOMIZE_REG_INIT
  wire  matchWay_prng_clock; // @[PRNG.scala 82:22]
  wire  matchWay_prng_reset; // @[PRNG.scala 82:22]
  wire  matchWay_prng_io_out_0; // @[PRNG.scala 82:22]
  wire  matchWay_prng_io_out_1; // @[PRNG.scala 82:22]
  wire  matchWay_prng_io_out_2; // @[PRNG.scala 82:22]
  reg [21:0] tag_0_0; // @[icache.scala 69:26]
  reg [21:0] tag_0_1; // @[icache.scala 69:26]
  reg [21:0] tag_0_2; // @[icache.scala 69:26]
  reg [21:0] tag_0_3; // @[icache.scala 69:26]
  reg [21:0] tag_0_4; // @[icache.scala 69:26]
  reg [21:0] tag_0_5; // @[icache.scala 69:26]
  reg [21:0] tag_0_6; // @[icache.scala 69:26]
  reg [21:0] tag_0_7; // @[icache.scala 69:26]
  reg [21:0] tag_0_8; // @[icache.scala 69:26]
  reg [21:0] tag_0_9; // @[icache.scala 69:26]
  reg [21:0] tag_0_10; // @[icache.scala 69:26]
  reg [21:0] tag_0_11; // @[icache.scala 69:26]
  reg [21:0] tag_0_12; // @[icache.scala 69:26]
  reg [21:0] tag_0_13; // @[icache.scala 69:26]
  reg [21:0] tag_0_14; // @[icache.scala 69:26]
  reg [21:0] tag_0_15; // @[icache.scala 69:26]
  reg [21:0] tag_1_0; // @[icache.scala 69:26]
  reg [21:0] tag_1_1; // @[icache.scala 69:26]
  reg [21:0] tag_1_2; // @[icache.scala 69:26]
  reg [21:0] tag_1_3; // @[icache.scala 69:26]
  reg [21:0] tag_1_4; // @[icache.scala 69:26]
  reg [21:0] tag_1_5; // @[icache.scala 69:26]
  reg [21:0] tag_1_6; // @[icache.scala 69:26]
  reg [21:0] tag_1_7; // @[icache.scala 69:26]
  reg [21:0] tag_1_8; // @[icache.scala 69:26]
  reg [21:0] tag_1_9; // @[icache.scala 69:26]
  reg [21:0] tag_1_10; // @[icache.scala 69:26]
  reg [21:0] tag_1_11; // @[icache.scala 69:26]
  reg [21:0] tag_1_12; // @[icache.scala 69:26]
  reg [21:0] tag_1_13; // @[icache.scala 69:26]
  reg [21:0] tag_1_14; // @[icache.scala 69:26]
  reg [21:0] tag_1_15; // @[icache.scala 69:26]
  reg [21:0] tag_2_0; // @[icache.scala 69:26]
  reg [21:0] tag_2_1; // @[icache.scala 69:26]
  reg [21:0] tag_2_2; // @[icache.scala 69:26]
  reg [21:0] tag_2_3; // @[icache.scala 69:26]
  reg [21:0] tag_2_4; // @[icache.scala 69:26]
  reg [21:0] tag_2_5; // @[icache.scala 69:26]
  reg [21:0] tag_2_6; // @[icache.scala 69:26]
  reg [21:0] tag_2_7; // @[icache.scala 69:26]
  reg [21:0] tag_2_8; // @[icache.scala 69:26]
  reg [21:0] tag_2_9; // @[icache.scala 69:26]
  reg [21:0] tag_2_10; // @[icache.scala 69:26]
  reg [21:0] tag_2_11; // @[icache.scala 69:26]
  reg [21:0] tag_2_12; // @[icache.scala 69:26]
  reg [21:0] tag_2_13; // @[icache.scala 69:26]
  reg [21:0] tag_2_14; // @[icache.scala 69:26]
  reg [21:0] tag_2_15; // @[icache.scala 69:26]
  reg [21:0] tag_3_0; // @[icache.scala 69:26]
  reg [21:0] tag_3_1; // @[icache.scala 69:26]
  reg [21:0] tag_3_2; // @[icache.scala 69:26]
  reg [21:0] tag_3_3; // @[icache.scala 69:26]
  reg [21:0] tag_3_4; // @[icache.scala 69:26]
  reg [21:0] tag_3_5; // @[icache.scala 69:26]
  reg [21:0] tag_3_6; // @[icache.scala 69:26]
  reg [21:0] tag_3_7; // @[icache.scala 69:26]
  reg [21:0] tag_3_8; // @[icache.scala 69:26]
  reg [21:0] tag_3_9; // @[icache.scala 69:26]
  reg [21:0] tag_3_10; // @[icache.scala 69:26]
  reg [21:0] tag_3_11; // @[icache.scala 69:26]
  reg [21:0] tag_3_12; // @[icache.scala 69:26]
  reg [21:0] tag_3_13; // @[icache.scala 69:26]
  reg [21:0] tag_3_14; // @[icache.scala 69:26]
  reg [21:0] tag_3_15; // @[icache.scala 69:26]
  reg  valid_0_0; // @[icache.scala 70:26]
  reg  valid_0_1; // @[icache.scala 70:26]
  reg  valid_0_2; // @[icache.scala 70:26]
  reg  valid_0_3; // @[icache.scala 70:26]
  reg  valid_0_4; // @[icache.scala 70:26]
  reg  valid_0_5; // @[icache.scala 70:26]
  reg  valid_0_6; // @[icache.scala 70:26]
  reg  valid_0_7; // @[icache.scala 70:26]
  reg  valid_0_8; // @[icache.scala 70:26]
  reg  valid_0_9; // @[icache.scala 70:26]
  reg  valid_0_10; // @[icache.scala 70:26]
  reg  valid_0_11; // @[icache.scala 70:26]
  reg  valid_0_12; // @[icache.scala 70:26]
  reg  valid_0_13; // @[icache.scala 70:26]
  reg  valid_0_14; // @[icache.scala 70:26]
  reg  valid_0_15; // @[icache.scala 70:26]
  reg  valid_1_0; // @[icache.scala 70:26]
  reg  valid_1_1; // @[icache.scala 70:26]
  reg  valid_1_2; // @[icache.scala 70:26]
  reg  valid_1_3; // @[icache.scala 70:26]
  reg  valid_1_4; // @[icache.scala 70:26]
  reg  valid_1_5; // @[icache.scala 70:26]
  reg  valid_1_6; // @[icache.scala 70:26]
  reg  valid_1_7; // @[icache.scala 70:26]
  reg  valid_1_8; // @[icache.scala 70:26]
  reg  valid_1_9; // @[icache.scala 70:26]
  reg  valid_1_10; // @[icache.scala 70:26]
  reg  valid_1_11; // @[icache.scala 70:26]
  reg  valid_1_12; // @[icache.scala 70:26]
  reg  valid_1_13; // @[icache.scala 70:26]
  reg  valid_1_14; // @[icache.scala 70:26]
  reg  valid_1_15; // @[icache.scala 70:26]
  reg  valid_2_0; // @[icache.scala 70:26]
  reg  valid_2_1; // @[icache.scala 70:26]
  reg  valid_2_2; // @[icache.scala 70:26]
  reg  valid_2_3; // @[icache.scala 70:26]
  reg  valid_2_4; // @[icache.scala 70:26]
  reg  valid_2_5; // @[icache.scala 70:26]
  reg  valid_2_6; // @[icache.scala 70:26]
  reg  valid_2_7; // @[icache.scala 70:26]
  reg  valid_2_8; // @[icache.scala 70:26]
  reg  valid_2_9; // @[icache.scala 70:26]
  reg  valid_2_10; // @[icache.scala 70:26]
  reg  valid_2_11; // @[icache.scala 70:26]
  reg  valid_2_12; // @[icache.scala 70:26]
  reg  valid_2_13; // @[icache.scala 70:26]
  reg  valid_2_14; // @[icache.scala 70:26]
  reg  valid_2_15; // @[icache.scala 70:26]
  reg  valid_3_0; // @[icache.scala 70:26]
  reg  valid_3_1; // @[icache.scala 70:26]
  reg  valid_3_2; // @[icache.scala 70:26]
  reg  valid_3_3; // @[icache.scala 70:26]
  reg  valid_3_4; // @[icache.scala 70:26]
  reg  valid_3_5; // @[icache.scala 70:26]
  reg  valid_3_6; // @[icache.scala 70:26]
  reg  valid_3_7; // @[icache.scala 70:26]
  reg  valid_3_8; // @[icache.scala 70:26]
  reg  valid_3_9; // @[icache.scala 70:26]
  reg  valid_3_10; // @[icache.scala 70:26]
  reg  valid_3_11; // @[icache.scala 70:26]
  reg  valid_3_12; // @[icache.scala 70:26]
  reg  valid_3_13; // @[icache.scala 70:26]
  reg  valid_3_14; // @[icache.scala 70:26]
  reg  valid_3_15; // @[icache.scala 70:26]
  reg  wait_r; // @[icache.scala 72:30]
  reg  valid_r; // @[icache.scala 73:30]
  wire  valid_in = io_icRead_arvalid & ~io_flush; // @[icache.scala 75:41]
  wire  hs_in = io_icRead_ready & io_icRead_arvalid; // @[icache.scala 76:39]
  wire  _io_icRead_ready_T = ~wait_r; // @[icache.scala 77:40]
  reg [31:0] addr_r; // @[icache.scala 79:34]
  reg [31:0] matchWay_r; // @[icache.scala 80:34]
  reg [2:0] axiOffset; // @[icache.scala 81:34]
  reg [63:0] databuf; // @[icache.scala 82:34]
  wire [31:0] cur_addr = hs_in ? io_icRead_addr : addr_r; // @[icache.scala 83:30]
  wire [21:0] instTag = cur_addr[31:10]; // @[icache.scala 84:35]
  wire [3:0] blockIdx = cur_addr[9:6]; // @[icache.scala 85:35]
  wire [5:0] cur_ram_addr = cur_addr[9:4]; // @[icache.scala 86:35]
  wire [1:0] cur_raddr_lo = axiOffset[2:1]; // @[icache.scala 87:100]
  wire [5:0] cur_raddr = {blockIdx,cur_raddr_lo}; // @[Cat.scala 30:58]
  wire [21:0] _GEN_1 = 4'h1 == blockIdx ? tag_0_1 : tag_0_0; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_2 = 4'h2 == blockIdx ? tag_0_2 : _GEN_1; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_3 = 4'h3 == blockIdx ? tag_0_3 : _GEN_2; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_4 = 4'h4 == blockIdx ? tag_0_4 : _GEN_3; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_5 = 4'h5 == blockIdx ? tag_0_5 : _GEN_4; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_6 = 4'h6 == blockIdx ? tag_0_6 : _GEN_5; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_7 = 4'h7 == blockIdx ? tag_0_7 : _GEN_6; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_8 = 4'h8 == blockIdx ? tag_0_8 : _GEN_7; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_9 = 4'h9 == blockIdx ? tag_0_9 : _GEN_8; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_10 = 4'ha == blockIdx ? tag_0_10 : _GEN_9; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_11 = 4'hb == blockIdx ? tag_0_11 : _GEN_10; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_12 = 4'hc == blockIdx ? tag_0_12 : _GEN_11; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_13 = 4'hd == blockIdx ? tag_0_13 : _GEN_12; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_14 = 4'he == blockIdx ? tag_0_14 : _GEN_13; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_15 = 4'hf == blockIdx ? tag_0_15 : _GEN_14; // @[icache.scala 88:85 icache.scala 88:85]
  wire  _GEN_17 = 4'h1 == blockIdx ? valid_0_1 : valid_0_0; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_18 = 4'h2 == blockIdx ? valid_0_2 : _GEN_17; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_19 = 4'h3 == blockIdx ? valid_0_3 : _GEN_18; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_20 = 4'h4 == blockIdx ? valid_0_4 : _GEN_19; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_21 = 4'h5 == blockIdx ? valid_0_5 : _GEN_20; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_22 = 4'h6 == blockIdx ? valid_0_6 : _GEN_21; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_23 = 4'h7 == blockIdx ? valid_0_7 : _GEN_22; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_24 = 4'h8 == blockIdx ? valid_0_8 : _GEN_23; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_25 = 4'h9 == blockIdx ? valid_0_9 : _GEN_24; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_26 = 4'ha == blockIdx ? valid_0_10 : _GEN_25; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_27 = 4'hb == blockIdx ? valid_0_11 : _GEN_26; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_28 = 4'hc == blockIdx ? valid_0_12 : _GEN_27; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_29 = 4'hd == blockIdx ? valid_0_13 : _GEN_28; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_30 = 4'he == blockIdx ? valid_0_14 : _GEN_29; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_31 = 4'hf == blockIdx ? valid_0_15 : _GEN_30; // @[icache.scala 88:97 icache.scala 88:97]
  wire  cache_hit_vec_0 = _GEN_15 == instTag & _GEN_31; // @[icache.scala 88:97]
  wire [21:0] _GEN_33 = 4'h1 == blockIdx ? tag_1_1 : tag_1_0; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_34 = 4'h2 == blockIdx ? tag_1_2 : _GEN_33; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_35 = 4'h3 == blockIdx ? tag_1_3 : _GEN_34; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_36 = 4'h4 == blockIdx ? tag_1_4 : _GEN_35; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_37 = 4'h5 == blockIdx ? tag_1_5 : _GEN_36; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_38 = 4'h6 == blockIdx ? tag_1_6 : _GEN_37; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_39 = 4'h7 == blockIdx ? tag_1_7 : _GEN_38; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_40 = 4'h8 == blockIdx ? tag_1_8 : _GEN_39; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_41 = 4'h9 == blockIdx ? tag_1_9 : _GEN_40; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_42 = 4'ha == blockIdx ? tag_1_10 : _GEN_41; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_43 = 4'hb == blockIdx ? tag_1_11 : _GEN_42; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_44 = 4'hc == blockIdx ? tag_1_12 : _GEN_43; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_45 = 4'hd == blockIdx ? tag_1_13 : _GEN_44; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_46 = 4'he == blockIdx ? tag_1_14 : _GEN_45; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_47 = 4'hf == blockIdx ? tag_1_15 : _GEN_46; // @[icache.scala 88:85 icache.scala 88:85]
  wire  _GEN_49 = 4'h1 == blockIdx ? valid_1_1 : valid_1_0; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_50 = 4'h2 == blockIdx ? valid_1_2 : _GEN_49; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_51 = 4'h3 == blockIdx ? valid_1_3 : _GEN_50; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_52 = 4'h4 == blockIdx ? valid_1_4 : _GEN_51; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_53 = 4'h5 == blockIdx ? valid_1_5 : _GEN_52; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_54 = 4'h6 == blockIdx ? valid_1_6 : _GEN_53; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_55 = 4'h7 == blockIdx ? valid_1_7 : _GEN_54; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_56 = 4'h8 == blockIdx ? valid_1_8 : _GEN_55; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_57 = 4'h9 == blockIdx ? valid_1_9 : _GEN_56; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_58 = 4'ha == blockIdx ? valid_1_10 : _GEN_57; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_59 = 4'hb == blockIdx ? valid_1_11 : _GEN_58; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_60 = 4'hc == blockIdx ? valid_1_12 : _GEN_59; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_61 = 4'hd == blockIdx ? valid_1_13 : _GEN_60; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_62 = 4'he == blockIdx ? valid_1_14 : _GEN_61; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_63 = 4'hf == blockIdx ? valid_1_15 : _GEN_62; // @[icache.scala 88:97 icache.scala 88:97]
  wire  cache_hit_vec_1 = _GEN_47 == instTag & _GEN_63; // @[icache.scala 88:97]
  wire [21:0] _GEN_65 = 4'h1 == blockIdx ? tag_2_1 : tag_2_0; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_66 = 4'h2 == blockIdx ? tag_2_2 : _GEN_65; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_67 = 4'h3 == blockIdx ? tag_2_3 : _GEN_66; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_68 = 4'h4 == blockIdx ? tag_2_4 : _GEN_67; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_69 = 4'h5 == blockIdx ? tag_2_5 : _GEN_68; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_70 = 4'h6 == blockIdx ? tag_2_6 : _GEN_69; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_71 = 4'h7 == blockIdx ? tag_2_7 : _GEN_70; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_72 = 4'h8 == blockIdx ? tag_2_8 : _GEN_71; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_73 = 4'h9 == blockIdx ? tag_2_9 : _GEN_72; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_74 = 4'ha == blockIdx ? tag_2_10 : _GEN_73; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_75 = 4'hb == blockIdx ? tag_2_11 : _GEN_74; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_76 = 4'hc == blockIdx ? tag_2_12 : _GEN_75; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_77 = 4'hd == blockIdx ? tag_2_13 : _GEN_76; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_78 = 4'he == blockIdx ? tag_2_14 : _GEN_77; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_79 = 4'hf == blockIdx ? tag_2_15 : _GEN_78; // @[icache.scala 88:85 icache.scala 88:85]
  wire  _GEN_81 = 4'h1 == blockIdx ? valid_2_1 : valid_2_0; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_82 = 4'h2 == blockIdx ? valid_2_2 : _GEN_81; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_83 = 4'h3 == blockIdx ? valid_2_3 : _GEN_82; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_84 = 4'h4 == blockIdx ? valid_2_4 : _GEN_83; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_85 = 4'h5 == blockIdx ? valid_2_5 : _GEN_84; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_86 = 4'h6 == blockIdx ? valid_2_6 : _GEN_85; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_87 = 4'h7 == blockIdx ? valid_2_7 : _GEN_86; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_88 = 4'h8 == blockIdx ? valid_2_8 : _GEN_87; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_89 = 4'h9 == blockIdx ? valid_2_9 : _GEN_88; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_90 = 4'ha == blockIdx ? valid_2_10 : _GEN_89; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_91 = 4'hb == blockIdx ? valid_2_11 : _GEN_90; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_92 = 4'hc == blockIdx ? valid_2_12 : _GEN_91; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_93 = 4'hd == blockIdx ? valid_2_13 : _GEN_92; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_94 = 4'he == blockIdx ? valid_2_14 : _GEN_93; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_95 = 4'hf == blockIdx ? valid_2_15 : _GEN_94; // @[icache.scala 88:97 icache.scala 88:97]
  wire  cache_hit_vec_2 = _GEN_79 == instTag & _GEN_95; // @[icache.scala 88:97]
  wire [21:0] _GEN_97 = 4'h1 == blockIdx ? tag_3_1 : tag_3_0; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_98 = 4'h2 == blockIdx ? tag_3_2 : _GEN_97; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_99 = 4'h3 == blockIdx ? tag_3_3 : _GEN_98; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_100 = 4'h4 == blockIdx ? tag_3_4 : _GEN_99; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_101 = 4'h5 == blockIdx ? tag_3_5 : _GEN_100; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_102 = 4'h6 == blockIdx ? tag_3_6 : _GEN_101; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_103 = 4'h7 == blockIdx ? tag_3_7 : _GEN_102; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_104 = 4'h8 == blockIdx ? tag_3_8 : _GEN_103; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_105 = 4'h9 == blockIdx ? tag_3_9 : _GEN_104; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_106 = 4'ha == blockIdx ? tag_3_10 : _GEN_105; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_107 = 4'hb == blockIdx ? tag_3_11 : _GEN_106; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_108 = 4'hc == blockIdx ? tag_3_12 : _GEN_107; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_109 = 4'hd == blockIdx ? tag_3_13 : _GEN_108; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_110 = 4'he == blockIdx ? tag_3_14 : _GEN_109; // @[icache.scala 88:85 icache.scala 88:85]
  wire [21:0] _GEN_111 = 4'hf == blockIdx ? tag_3_15 : _GEN_110; // @[icache.scala 88:85 icache.scala 88:85]
  wire  _GEN_113 = 4'h1 == blockIdx ? valid_3_1 : valid_3_0; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_114 = 4'h2 == blockIdx ? valid_3_2 : _GEN_113; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_115 = 4'h3 == blockIdx ? valid_3_3 : _GEN_114; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_116 = 4'h4 == blockIdx ? valid_3_4 : _GEN_115; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_117 = 4'h5 == blockIdx ? valid_3_5 : _GEN_116; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_118 = 4'h6 == blockIdx ? valid_3_6 : _GEN_117; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_119 = 4'h7 == blockIdx ? valid_3_7 : _GEN_118; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_120 = 4'h8 == blockIdx ? valid_3_8 : _GEN_119; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_121 = 4'h9 == blockIdx ? valid_3_9 : _GEN_120; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_122 = 4'ha == blockIdx ? valid_3_10 : _GEN_121; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_123 = 4'hb == blockIdx ? valid_3_11 : _GEN_122; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_124 = 4'hc == blockIdx ? valid_3_12 : _GEN_123; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_125 = 4'hd == blockIdx ? valid_3_13 : _GEN_124; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_126 = 4'he == blockIdx ? valid_3_14 : _GEN_125; // @[icache.scala 88:97 icache.scala 88:97]
  wire  _GEN_127 = 4'hf == blockIdx ? valid_3_15 : _GEN_126; // @[icache.scala 88:97 icache.scala 88:97]
  wire  cache_hit_vec_3 = _GEN_111 == instTag & _GEN_127; // @[icache.scala 88:97]
  wire [3:0] _cacheHit_T = {cache_hit_vec_3,cache_hit_vec_2,cache_hit_vec_1,cache_hit_vec_0}; // @[icache.scala 89:47]
  wire  cacheHit = |_cacheHit_T; // @[icache.scala 89:50]
  wire [1:0] matchWay_hi_1 = _cacheHit_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] matchWay_lo_1 = _cacheHit_T[1:0]; // @[OneHot.scala 31:18]
  wire  matchWay_hi_2 = |matchWay_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _matchWay_T_1 = matchWay_hi_1 | matchWay_lo_1; // @[OneHot.scala 32:28]
  wire  matchWay_lo_2 = _matchWay_T_1[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] _matchWay_T_2 = {matchWay_hi_2,matchWay_lo_2}; // @[Cat.scala 30:58]
  wire [2:0] _matchWay_T_3 = {matchWay_prng_io_out_2,matchWay_prng_io_out_1,matchWay_prng_io_out_0}; // @[PRNG.scala 86:17]
  wire [1:0] matchWay = cacheHit ? _matchWay_T_2 : _matchWay_T_3[2:1]; // @[icache.scala 90:30]
  wire [31:0] cur_way = hs_in ? {{30'd0}, matchWay} : matchWay_r; // @[icache.scala 91:30]
  wire [3:0] pre_blockIdx = addr_r[9:6]; // @[icache.scala 92:33]
  wire [21:0] pre_instTag = addr_r[31:10]; // @[icache.scala 93:33]
  wire  _GEN_130 = io_flush ? 1'h0 : valid_0_0; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_131 = io_flush ? 1'h0 : valid_0_1; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_132 = io_flush ? 1'h0 : valid_0_2; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_133 = io_flush ? 1'h0 : valid_0_3; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_134 = io_flush ? 1'h0 : valid_0_4; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_135 = io_flush ? 1'h0 : valid_0_5; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_136 = io_flush ? 1'h0 : valid_0_6; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_137 = io_flush ? 1'h0 : valid_0_7; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_138 = io_flush ? 1'h0 : valid_0_8; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_139 = io_flush ? 1'h0 : valid_0_9; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_140 = io_flush ? 1'h0 : valid_0_10; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_141 = io_flush ? 1'h0 : valid_0_11; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_142 = io_flush ? 1'h0 : valid_0_12; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_143 = io_flush ? 1'h0 : valid_0_13; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_144 = io_flush ? 1'h0 : valid_0_14; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_145 = io_flush ? 1'h0 : valid_0_15; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_146 = io_flush ? 1'h0 : valid_1_0; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_147 = io_flush ? 1'h0 : valid_1_1; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_148 = io_flush ? 1'h0 : valid_1_2; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_149 = io_flush ? 1'h0 : valid_1_3; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_150 = io_flush ? 1'h0 : valid_1_4; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_151 = io_flush ? 1'h0 : valid_1_5; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_152 = io_flush ? 1'h0 : valid_1_6; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_153 = io_flush ? 1'h0 : valid_1_7; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_154 = io_flush ? 1'h0 : valid_1_8; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_155 = io_flush ? 1'h0 : valid_1_9; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_156 = io_flush ? 1'h0 : valid_1_10; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_157 = io_flush ? 1'h0 : valid_1_11; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_158 = io_flush ? 1'h0 : valid_1_12; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_159 = io_flush ? 1'h0 : valid_1_13; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_160 = io_flush ? 1'h0 : valid_1_14; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_161 = io_flush ? 1'h0 : valid_1_15; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_162 = io_flush ? 1'h0 : valid_2_0; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_163 = io_flush ? 1'h0 : valid_2_1; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_164 = io_flush ? 1'h0 : valid_2_2; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_165 = io_flush ? 1'h0 : valid_2_3; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_166 = io_flush ? 1'h0 : valid_2_4; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_167 = io_flush ? 1'h0 : valid_2_5; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_168 = io_flush ? 1'h0 : valid_2_6; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_169 = io_flush ? 1'h0 : valid_2_7; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_170 = io_flush ? 1'h0 : valid_2_8; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_171 = io_flush ? 1'h0 : valid_2_9; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_172 = io_flush ? 1'h0 : valid_2_10; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_173 = io_flush ? 1'h0 : valid_2_11; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_174 = io_flush ? 1'h0 : valid_2_12; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_175 = io_flush ? 1'h0 : valid_2_13; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_176 = io_flush ? 1'h0 : valid_2_14; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_177 = io_flush ? 1'h0 : valid_2_15; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_178 = io_flush ? 1'h0 : valid_3_0; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_179 = io_flush ? 1'h0 : valid_3_1; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_180 = io_flush ? 1'h0 : valid_3_2; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_181 = io_flush ? 1'h0 : valid_3_3; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_182 = io_flush ? 1'h0 : valid_3_4; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_183 = io_flush ? 1'h0 : valid_3_5; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_184 = io_flush ? 1'h0 : valid_3_6; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_185 = io_flush ? 1'h0 : valid_3_7; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_186 = io_flush ? 1'h0 : valid_3_8; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_187 = io_flush ? 1'h0 : valid_3_9; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_188 = io_flush ? 1'h0 : valid_3_10; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_189 = io_flush ? 1'h0 : valid_3_11; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_190 = io_flush ? 1'h0 : valid_3_12; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_191 = io_flush ? 1'h0 : valid_3_13; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_192 = io_flush ? 1'h0 : valid_3_14; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  wire  _GEN_193 = io_flush ? 1'h0 : valid_3_15; // @[icache.scala 99:19 icache.scala 100:17 icache.scala 70:26]
  reg [1:0] state; // @[icache.scala 103:24]
  wire [127:0] _rdata128_T_1 = 32'h0 == matchWay_r ? io_ic2sr0_rdata : 128'h0; // @[Mux.scala 80:57]
  wire [127:0] _rdata128_T_3 = 32'h1 == matchWay_r ? io_ic2sr1_rdata : _rdata128_T_1; // @[Mux.scala 80:57]
  wire [127:0] _rdata128_T_5 = 32'h2 == matchWay_r ? io_ic2sr2_rdata : _rdata128_T_3; // @[Mux.scala 80:57]
  wire [127:0] rdata128 = 32'h3 == matchWay_r ? io_ic2sr3_rdata : _rdata128_T_5; // @[Mux.scala 80:57]
  wire  _io_ic2sr0_cen_T_1 = wait_r | hs_in; // @[icache.scala 120:52]
  wire  _T = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_6 = 2'h2 == state; // @[Conditional.scala 37:30]
  reg  rdataEn; // @[icache.scala 140:30]
  wire  _GEN_470 = rdataEn & io_instAxi_rd_valid & axiOffset[0]; // @[icache.scala 166:49 icache.scala 136:13]
  wire  _GEN_739 = _T_4 ? 1'h0 : _T_6 & _GEN_470; // @[Conditional.scala 39:67 icache.scala 136:13]
  wire  wen = _T ? 1'h0 : _GEN_739; // @[Conditional.scala 40:58 icache.scala 136:13]
  reg  raddrEn; // @[icache.scala 138:30]
  reg [31:0] raddr; // @[icache.scala 139:30]
  wire [31:0] _raddr_T = cur_addr & 32'hffffffc0; // @[icache.scala 150:37]
  wire  _GEN_199 = ~hs_in & _io_icRead_ready_T ? 1'h0 : cacheHit; // @[icache.scala 144:36 icache.scala 74:13]
  wire  _GEN_206 = raddrEn & io_instAxi_ra_ready | rdataEn; // @[icache.scala 158:49 icache.scala 161:25 icache.scala 140:30]
  wire [2:0] _axiOffset_T_1 = axiOffset + 3'h1; // @[icache.scala 167:40]
  wire [63:0] _GEN_209 = axiOffset[0] ? databuf : io_instAxi_rd_bits_data; // @[icache.scala 168:35 icache.scala 82:34 icache.scala 171:29]
  wire  _GEN_1006 = 2'h0 == matchWay_r[1:0]; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1007 = 4'h0 == pre_blockIdx; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_210 = 2'h0 == matchWay_r[1:0] & 4'h0 == pre_blockIdx ? pre_instTag : tag_0_0; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1009 = 4'h1 == pre_blockIdx; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_211 = 2'h0 == matchWay_r[1:0] & 4'h1 == pre_blockIdx ? pre_instTag : tag_0_1; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1011 = 4'h2 == pre_blockIdx; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_212 = 2'h0 == matchWay_r[1:0] & 4'h2 == pre_blockIdx ? pre_instTag : tag_0_2; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1013 = 4'h3 == pre_blockIdx; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_213 = 2'h0 == matchWay_r[1:0] & 4'h3 == pre_blockIdx ? pre_instTag : tag_0_3; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1015 = 4'h4 == pre_blockIdx; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_214 = 2'h0 == matchWay_r[1:0] & 4'h4 == pre_blockIdx ? pre_instTag : tag_0_4; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1017 = 4'h5 == pre_blockIdx; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_215 = 2'h0 == matchWay_r[1:0] & 4'h5 == pre_blockIdx ? pre_instTag : tag_0_5; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1019 = 4'h6 == pre_blockIdx; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_216 = 2'h0 == matchWay_r[1:0] & 4'h6 == pre_blockIdx ? pre_instTag : tag_0_6; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1021 = 4'h7 == pre_blockIdx; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_217 = 2'h0 == matchWay_r[1:0] & 4'h7 == pre_blockIdx ? pre_instTag : tag_0_7; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1023 = 4'h8 == pre_blockIdx; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_218 = 2'h0 == matchWay_r[1:0] & 4'h8 == pre_blockIdx ? pre_instTag : tag_0_8; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1025 = 4'h9 == pre_blockIdx; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_219 = 2'h0 == matchWay_r[1:0] & 4'h9 == pre_blockIdx ? pre_instTag : tag_0_9; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1027 = 4'ha == pre_blockIdx; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_220 = 2'h0 == matchWay_r[1:0] & 4'ha == pre_blockIdx ? pre_instTag : tag_0_10; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1029 = 4'hb == pre_blockIdx; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_221 = 2'h0 == matchWay_r[1:0] & 4'hb == pre_blockIdx ? pre_instTag : tag_0_11; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1031 = 4'hc == pre_blockIdx; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_222 = 2'h0 == matchWay_r[1:0] & 4'hc == pre_blockIdx ? pre_instTag : tag_0_12; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1033 = 4'hd == pre_blockIdx; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_223 = 2'h0 == matchWay_r[1:0] & 4'hd == pre_blockIdx ? pre_instTag : tag_0_13; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1035 = 4'he == pre_blockIdx; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_224 = 2'h0 == matchWay_r[1:0] & 4'he == pre_blockIdx ? pre_instTag : tag_0_14; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1037 = 4'hf == pre_blockIdx; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_225 = 2'h0 == matchWay_r[1:0] & 4'hf == pre_blockIdx ? pre_instTag : tag_0_15; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1038 = 2'h1 == matchWay_r[1:0]; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_226 = 2'h1 == matchWay_r[1:0] & 4'h0 == pre_blockIdx ? pre_instTag : tag_1_0; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_227 = 2'h1 == matchWay_r[1:0] & 4'h1 == pre_blockIdx ? pre_instTag : tag_1_1; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_228 = 2'h1 == matchWay_r[1:0] & 4'h2 == pre_blockIdx ? pre_instTag : tag_1_2; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_229 = 2'h1 == matchWay_r[1:0] & 4'h3 == pre_blockIdx ? pre_instTag : tag_1_3; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_230 = 2'h1 == matchWay_r[1:0] & 4'h4 == pre_blockIdx ? pre_instTag : tag_1_4; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_231 = 2'h1 == matchWay_r[1:0] & 4'h5 == pre_blockIdx ? pre_instTag : tag_1_5; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_232 = 2'h1 == matchWay_r[1:0] & 4'h6 == pre_blockIdx ? pre_instTag : tag_1_6; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_233 = 2'h1 == matchWay_r[1:0] & 4'h7 == pre_blockIdx ? pre_instTag : tag_1_7; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_234 = 2'h1 == matchWay_r[1:0] & 4'h8 == pre_blockIdx ? pre_instTag : tag_1_8; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_235 = 2'h1 == matchWay_r[1:0] & 4'h9 == pre_blockIdx ? pre_instTag : tag_1_9; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_236 = 2'h1 == matchWay_r[1:0] & 4'ha == pre_blockIdx ? pre_instTag : tag_1_10; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_237 = 2'h1 == matchWay_r[1:0] & 4'hb == pre_blockIdx ? pre_instTag : tag_1_11; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_238 = 2'h1 == matchWay_r[1:0] & 4'hc == pre_blockIdx ? pre_instTag : tag_1_12; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_239 = 2'h1 == matchWay_r[1:0] & 4'hd == pre_blockIdx ? pre_instTag : tag_1_13; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_240 = 2'h1 == matchWay_r[1:0] & 4'he == pre_blockIdx ? pre_instTag : tag_1_14; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_241 = 2'h1 == matchWay_r[1:0] & 4'hf == pre_blockIdx ? pre_instTag : tag_1_15; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1070 = 2'h2 == matchWay_r[1:0]; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_242 = 2'h2 == matchWay_r[1:0] & 4'h0 == pre_blockIdx ? pre_instTag : tag_2_0; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_243 = 2'h2 == matchWay_r[1:0] & 4'h1 == pre_blockIdx ? pre_instTag : tag_2_1; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_244 = 2'h2 == matchWay_r[1:0] & 4'h2 == pre_blockIdx ? pre_instTag : tag_2_2; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_245 = 2'h2 == matchWay_r[1:0] & 4'h3 == pre_blockIdx ? pre_instTag : tag_2_3; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_246 = 2'h2 == matchWay_r[1:0] & 4'h4 == pre_blockIdx ? pre_instTag : tag_2_4; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_247 = 2'h2 == matchWay_r[1:0] & 4'h5 == pre_blockIdx ? pre_instTag : tag_2_5; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_248 = 2'h2 == matchWay_r[1:0] & 4'h6 == pre_blockIdx ? pre_instTag : tag_2_6; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_249 = 2'h2 == matchWay_r[1:0] & 4'h7 == pre_blockIdx ? pre_instTag : tag_2_7; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_250 = 2'h2 == matchWay_r[1:0] & 4'h8 == pre_blockIdx ? pre_instTag : tag_2_8; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_251 = 2'h2 == matchWay_r[1:0] & 4'h9 == pre_blockIdx ? pre_instTag : tag_2_9; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_252 = 2'h2 == matchWay_r[1:0] & 4'ha == pre_blockIdx ? pre_instTag : tag_2_10; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_253 = 2'h2 == matchWay_r[1:0] & 4'hb == pre_blockIdx ? pre_instTag : tag_2_11; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_254 = 2'h2 == matchWay_r[1:0] & 4'hc == pre_blockIdx ? pre_instTag : tag_2_12; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_255 = 2'h2 == matchWay_r[1:0] & 4'hd == pre_blockIdx ? pre_instTag : tag_2_13; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_256 = 2'h2 == matchWay_r[1:0] & 4'he == pre_blockIdx ? pre_instTag : tag_2_14; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_257 = 2'h2 == matchWay_r[1:0] & 4'hf == pre_blockIdx ? pre_instTag : tag_2_15; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_1102 = 2'h3 == matchWay_r[1:0]; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_258 = 2'h3 == matchWay_r[1:0] & 4'h0 == pre_blockIdx ? pre_instTag : tag_3_0; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_259 = 2'h3 == matchWay_r[1:0] & 4'h1 == pre_blockIdx ? pre_instTag : tag_3_1; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_260 = 2'h3 == matchWay_r[1:0] & 4'h2 == pre_blockIdx ? pre_instTag : tag_3_2; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_261 = 2'h3 == matchWay_r[1:0] & 4'h3 == pre_blockIdx ? pre_instTag : tag_3_3; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_262 = 2'h3 == matchWay_r[1:0] & 4'h4 == pre_blockIdx ? pre_instTag : tag_3_4; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_263 = 2'h3 == matchWay_r[1:0] & 4'h5 == pre_blockIdx ? pre_instTag : tag_3_5; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_264 = 2'h3 == matchWay_r[1:0] & 4'h6 == pre_blockIdx ? pre_instTag : tag_3_6; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_265 = 2'h3 == matchWay_r[1:0] & 4'h7 == pre_blockIdx ? pre_instTag : tag_3_7; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_266 = 2'h3 == matchWay_r[1:0] & 4'h8 == pre_blockIdx ? pre_instTag : tag_3_8; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_267 = 2'h3 == matchWay_r[1:0] & 4'h9 == pre_blockIdx ? pre_instTag : tag_3_9; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_268 = 2'h3 == matchWay_r[1:0] & 4'ha == pre_blockIdx ? pre_instTag : tag_3_10; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_269 = 2'h3 == matchWay_r[1:0] & 4'hb == pre_blockIdx ? pre_instTag : tag_3_11; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_270 = 2'h3 == matchWay_r[1:0] & 4'hc == pre_blockIdx ? pre_instTag : tag_3_12; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_271 = 2'h3 == matchWay_r[1:0] & 4'hd == pre_blockIdx ? pre_instTag : tag_3_13; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_272 = 2'h3 == matchWay_r[1:0] & 4'he == pre_blockIdx ? pre_instTag : tag_3_14; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire [21:0] _GEN_273 = 2'h3 == matchWay_r[1:0] & 4'hf == pre_blockIdx ? pre_instTag : tag_3_15; // @[icache.scala 175:51 icache.scala 175:51 icache.scala 69:26]
  wire  _GEN_274 = _GEN_1006 & _GEN_1007 | _GEN_130; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_275 = _GEN_1006 & _GEN_1009 | _GEN_131; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_276 = _GEN_1006 & _GEN_1011 | _GEN_132; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_277 = _GEN_1006 & _GEN_1013 | _GEN_133; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_278 = _GEN_1006 & _GEN_1015 | _GEN_134; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_279 = _GEN_1006 & _GEN_1017 | _GEN_135; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_280 = _GEN_1006 & _GEN_1019 | _GEN_136; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_281 = _GEN_1006 & _GEN_1021 | _GEN_137; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_282 = _GEN_1006 & _GEN_1023 | _GEN_138; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_283 = _GEN_1006 & _GEN_1025 | _GEN_139; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_284 = _GEN_1006 & _GEN_1027 | _GEN_140; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_285 = _GEN_1006 & _GEN_1029 | _GEN_141; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_286 = _GEN_1006 & _GEN_1031 | _GEN_142; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_287 = _GEN_1006 & _GEN_1033 | _GEN_143; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_288 = _GEN_1006 & _GEN_1035 | _GEN_144; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_289 = _GEN_1006 & _GEN_1037 | _GEN_145; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_290 = _GEN_1038 & _GEN_1007 | _GEN_146; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_291 = _GEN_1038 & _GEN_1009 | _GEN_147; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_292 = _GEN_1038 & _GEN_1011 | _GEN_148; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_293 = _GEN_1038 & _GEN_1013 | _GEN_149; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_294 = _GEN_1038 & _GEN_1015 | _GEN_150; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_295 = _GEN_1038 & _GEN_1017 | _GEN_151; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_296 = _GEN_1038 & _GEN_1019 | _GEN_152; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_297 = _GEN_1038 & _GEN_1021 | _GEN_153; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_298 = _GEN_1038 & _GEN_1023 | _GEN_154; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_299 = _GEN_1038 & _GEN_1025 | _GEN_155; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_300 = _GEN_1038 & _GEN_1027 | _GEN_156; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_301 = _GEN_1038 & _GEN_1029 | _GEN_157; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_302 = _GEN_1038 & _GEN_1031 | _GEN_158; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_303 = _GEN_1038 & _GEN_1033 | _GEN_159; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_304 = _GEN_1038 & _GEN_1035 | _GEN_160; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_305 = _GEN_1038 & _GEN_1037 | _GEN_161; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_306 = _GEN_1070 & _GEN_1007 | _GEN_162; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_307 = _GEN_1070 & _GEN_1009 | _GEN_163; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_308 = _GEN_1070 & _GEN_1011 | _GEN_164; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_309 = _GEN_1070 & _GEN_1013 | _GEN_165; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_310 = _GEN_1070 & _GEN_1015 | _GEN_166; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_311 = _GEN_1070 & _GEN_1017 | _GEN_167; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_312 = _GEN_1070 & _GEN_1019 | _GEN_168; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_313 = _GEN_1070 & _GEN_1021 | _GEN_169; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_314 = _GEN_1070 & _GEN_1023 | _GEN_170; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_315 = _GEN_1070 & _GEN_1025 | _GEN_171; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_316 = _GEN_1070 & _GEN_1027 | _GEN_172; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_317 = _GEN_1070 & _GEN_1029 | _GEN_173; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_318 = _GEN_1070 & _GEN_1031 | _GEN_174; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_319 = _GEN_1070 & _GEN_1033 | _GEN_175; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_320 = _GEN_1070 & _GEN_1035 | _GEN_176; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_321 = _GEN_1070 & _GEN_1037 | _GEN_177; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_322 = _GEN_1102 & _GEN_1007 | _GEN_178; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_323 = _GEN_1102 & _GEN_1009 | _GEN_179; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_324 = _GEN_1102 & _GEN_1011 | _GEN_180; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_325 = _GEN_1102 & _GEN_1013 | _GEN_181; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_326 = _GEN_1102 & _GEN_1015 | _GEN_182; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_327 = _GEN_1102 & _GEN_1017 | _GEN_183; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_328 = _GEN_1102 & _GEN_1019 | _GEN_184; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_329 = _GEN_1102 & _GEN_1021 | _GEN_185; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_330 = _GEN_1102 & _GEN_1023 | _GEN_186; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_331 = _GEN_1102 & _GEN_1025 | _GEN_187; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_332 = _GEN_1102 & _GEN_1027 | _GEN_188; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_333 = _GEN_1102 & _GEN_1029 | _GEN_189; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_334 = _GEN_1102 & _GEN_1031 | _GEN_190; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_335 = _GEN_1102 & _GEN_1033 | _GEN_191; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_336 = _GEN_1102 & _GEN_1035 | _GEN_192; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_337 = _GEN_1102 & _GEN_1037 | _GEN_193; // @[icache.scala 176:53 icache.scala 176:53]
  wire  _GEN_338 = io_instAxi_rd_bits_last ? 1'h0 : rdataEn; // @[icache.scala 173:46 icache.scala 174:29 icache.scala 140:30]
  wire [21:0] _GEN_339 = io_instAxi_rd_bits_last ? _GEN_210 : tag_0_0; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_340 = io_instAxi_rd_bits_last ? _GEN_211 : tag_0_1; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_341 = io_instAxi_rd_bits_last ? _GEN_212 : tag_0_2; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_342 = io_instAxi_rd_bits_last ? _GEN_213 : tag_0_3; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_343 = io_instAxi_rd_bits_last ? _GEN_214 : tag_0_4; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_344 = io_instAxi_rd_bits_last ? _GEN_215 : tag_0_5; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_345 = io_instAxi_rd_bits_last ? _GEN_216 : tag_0_6; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_346 = io_instAxi_rd_bits_last ? _GEN_217 : tag_0_7; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_347 = io_instAxi_rd_bits_last ? _GEN_218 : tag_0_8; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_348 = io_instAxi_rd_bits_last ? _GEN_219 : tag_0_9; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_349 = io_instAxi_rd_bits_last ? _GEN_220 : tag_0_10; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_350 = io_instAxi_rd_bits_last ? _GEN_221 : tag_0_11; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_351 = io_instAxi_rd_bits_last ? _GEN_222 : tag_0_12; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_352 = io_instAxi_rd_bits_last ? _GEN_223 : tag_0_13; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_353 = io_instAxi_rd_bits_last ? _GEN_224 : tag_0_14; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_354 = io_instAxi_rd_bits_last ? _GEN_225 : tag_0_15; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_355 = io_instAxi_rd_bits_last ? _GEN_226 : tag_1_0; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_356 = io_instAxi_rd_bits_last ? _GEN_227 : tag_1_1; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_357 = io_instAxi_rd_bits_last ? _GEN_228 : tag_1_2; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_358 = io_instAxi_rd_bits_last ? _GEN_229 : tag_1_3; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_359 = io_instAxi_rd_bits_last ? _GEN_230 : tag_1_4; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_360 = io_instAxi_rd_bits_last ? _GEN_231 : tag_1_5; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_361 = io_instAxi_rd_bits_last ? _GEN_232 : tag_1_6; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_362 = io_instAxi_rd_bits_last ? _GEN_233 : tag_1_7; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_363 = io_instAxi_rd_bits_last ? _GEN_234 : tag_1_8; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_364 = io_instAxi_rd_bits_last ? _GEN_235 : tag_1_9; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_365 = io_instAxi_rd_bits_last ? _GEN_236 : tag_1_10; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_366 = io_instAxi_rd_bits_last ? _GEN_237 : tag_1_11; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_367 = io_instAxi_rd_bits_last ? _GEN_238 : tag_1_12; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_368 = io_instAxi_rd_bits_last ? _GEN_239 : tag_1_13; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_369 = io_instAxi_rd_bits_last ? _GEN_240 : tag_1_14; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_370 = io_instAxi_rd_bits_last ? _GEN_241 : tag_1_15; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_371 = io_instAxi_rd_bits_last ? _GEN_242 : tag_2_0; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_372 = io_instAxi_rd_bits_last ? _GEN_243 : tag_2_1; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_373 = io_instAxi_rd_bits_last ? _GEN_244 : tag_2_2; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_374 = io_instAxi_rd_bits_last ? _GEN_245 : tag_2_3; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_375 = io_instAxi_rd_bits_last ? _GEN_246 : tag_2_4; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_376 = io_instAxi_rd_bits_last ? _GEN_247 : tag_2_5; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_377 = io_instAxi_rd_bits_last ? _GEN_248 : tag_2_6; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_378 = io_instAxi_rd_bits_last ? _GEN_249 : tag_2_7; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_379 = io_instAxi_rd_bits_last ? _GEN_250 : tag_2_8; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_380 = io_instAxi_rd_bits_last ? _GEN_251 : tag_2_9; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_381 = io_instAxi_rd_bits_last ? _GEN_252 : tag_2_10; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_382 = io_instAxi_rd_bits_last ? _GEN_253 : tag_2_11; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_383 = io_instAxi_rd_bits_last ? _GEN_254 : tag_2_12; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_384 = io_instAxi_rd_bits_last ? _GEN_255 : tag_2_13; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_385 = io_instAxi_rd_bits_last ? _GEN_256 : tag_2_14; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_386 = io_instAxi_rd_bits_last ? _GEN_257 : tag_2_15; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_387 = io_instAxi_rd_bits_last ? _GEN_258 : tag_3_0; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_388 = io_instAxi_rd_bits_last ? _GEN_259 : tag_3_1; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_389 = io_instAxi_rd_bits_last ? _GEN_260 : tag_3_2; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_390 = io_instAxi_rd_bits_last ? _GEN_261 : tag_3_3; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_391 = io_instAxi_rd_bits_last ? _GEN_262 : tag_3_4; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_392 = io_instAxi_rd_bits_last ? _GEN_263 : tag_3_5; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_393 = io_instAxi_rd_bits_last ? _GEN_264 : tag_3_6; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_394 = io_instAxi_rd_bits_last ? _GEN_265 : tag_3_7; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_395 = io_instAxi_rd_bits_last ? _GEN_266 : tag_3_8; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_396 = io_instAxi_rd_bits_last ? _GEN_267 : tag_3_9; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_397 = io_instAxi_rd_bits_last ? _GEN_268 : tag_3_10; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_398 = io_instAxi_rd_bits_last ? _GEN_269 : tag_3_11; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_399 = io_instAxi_rd_bits_last ? _GEN_270 : tag_3_12; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_400 = io_instAxi_rd_bits_last ? _GEN_271 : tag_3_13; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_401 = io_instAxi_rd_bits_last ? _GEN_272 : tag_3_14; // @[icache.scala 173:46 icache.scala 69:26]
  wire [21:0] _GEN_402 = io_instAxi_rd_bits_last ? _GEN_273 : tag_3_15; // @[icache.scala 173:46 icache.scala 69:26]
  wire  _GEN_403 = io_instAxi_rd_bits_last ? _GEN_274 : _GEN_130; // @[icache.scala 173:46]
  wire  _GEN_404 = io_instAxi_rd_bits_last ? _GEN_275 : _GEN_131; // @[icache.scala 173:46]
  wire  _GEN_405 = io_instAxi_rd_bits_last ? _GEN_276 : _GEN_132; // @[icache.scala 173:46]
  wire  _GEN_406 = io_instAxi_rd_bits_last ? _GEN_277 : _GEN_133; // @[icache.scala 173:46]
  wire  _GEN_407 = io_instAxi_rd_bits_last ? _GEN_278 : _GEN_134; // @[icache.scala 173:46]
  wire  _GEN_408 = io_instAxi_rd_bits_last ? _GEN_279 : _GEN_135; // @[icache.scala 173:46]
  wire  _GEN_409 = io_instAxi_rd_bits_last ? _GEN_280 : _GEN_136; // @[icache.scala 173:46]
  wire  _GEN_410 = io_instAxi_rd_bits_last ? _GEN_281 : _GEN_137; // @[icache.scala 173:46]
  wire  _GEN_411 = io_instAxi_rd_bits_last ? _GEN_282 : _GEN_138; // @[icache.scala 173:46]
  wire  _GEN_412 = io_instAxi_rd_bits_last ? _GEN_283 : _GEN_139; // @[icache.scala 173:46]
  wire  _GEN_413 = io_instAxi_rd_bits_last ? _GEN_284 : _GEN_140; // @[icache.scala 173:46]
  wire  _GEN_414 = io_instAxi_rd_bits_last ? _GEN_285 : _GEN_141; // @[icache.scala 173:46]
  wire  _GEN_415 = io_instAxi_rd_bits_last ? _GEN_286 : _GEN_142; // @[icache.scala 173:46]
  wire  _GEN_416 = io_instAxi_rd_bits_last ? _GEN_287 : _GEN_143; // @[icache.scala 173:46]
  wire  _GEN_417 = io_instAxi_rd_bits_last ? _GEN_288 : _GEN_144; // @[icache.scala 173:46]
  wire  _GEN_418 = io_instAxi_rd_bits_last ? _GEN_289 : _GEN_145; // @[icache.scala 173:46]
  wire  _GEN_419 = io_instAxi_rd_bits_last ? _GEN_290 : _GEN_146; // @[icache.scala 173:46]
  wire  _GEN_420 = io_instAxi_rd_bits_last ? _GEN_291 : _GEN_147; // @[icache.scala 173:46]
  wire  _GEN_421 = io_instAxi_rd_bits_last ? _GEN_292 : _GEN_148; // @[icache.scala 173:46]
  wire  _GEN_422 = io_instAxi_rd_bits_last ? _GEN_293 : _GEN_149; // @[icache.scala 173:46]
  wire  _GEN_423 = io_instAxi_rd_bits_last ? _GEN_294 : _GEN_150; // @[icache.scala 173:46]
  wire  _GEN_424 = io_instAxi_rd_bits_last ? _GEN_295 : _GEN_151; // @[icache.scala 173:46]
  wire  _GEN_425 = io_instAxi_rd_bits_last ? _GEN_296 : _GEN_152; // @[icache.scala 173:46]
  wire  _GEN_426 = io_instAxi_rd_bits_last ? _GEN_297 : _GEN_153; // @[icache.scala 173:46]
  wire  _GEN_427 = io_instAxi_rd_bits_last ? _GEN_298 : _GEN_154; // @[icache.scala 173:46]
  wire  _GEN_428 = io_instAxi_rd_bits_last ? _GEN_299 : _GEN_155; // @[icache.scala 173:46]
  wire  _GEN_429 = io_instAxi_rd_bits_last ? _GEN_300 : _GEN_156; // @[icache.scala 173:46]
  wire  _GEN_430 = io_instAxi_rd_bits_last ? _GEN_301 : _GEN_157; // @[icache.scala 173:46]
  wire  _GEN_431 = io_instAxi_rd_bits_last ? _GEN_302 : _GEN_158; // @[icache.scala 173:46]
  wire  _GEN_432 = io_instAxi_rd_bits_last ? _GEN_303 : _GEN_159; // @[icache.scala 173:46]
  wire  _GEN_433 = io_instAxi_rd_bits_last ? _GEN_304 : _GEN_160; // @[icache.scala 173:46]
  wire  _GEN_434 = io_instAxi_rd_bits_last ? _GEN_305 : _GEN_161; // @[icache.scala 173:46]
  wire  _GEN_435 = io_instAxi_rd_bits_last ? _GEN_306 : _GEN_162; // @[icache.scala 173:46]
  wire  _GEN_436 = io_instAxi_rd_bits_last ? _GEN_307 : _GEN_163; // @[icache.scala 173:46]
  wire  _GEN_437 = io_instAxi_rd_bits_last ? _GEN_308 : _GEN_164; // @[icache.scala 173:46]
  wire  _GEN_438 = io_instAxi_rd_bits_last ? _GEN_309 : _GEN_165; // @[icache.scala 173:46]
  wire  _GEN_439 = io_instAxi_rd_bits_last ? _GEN_310 : _GEN_166; // @[icache.scala 173:46]
  wire  _GEN_440 = io_instAxi_rd_bits_last ? _GEN_311 : _GEN_167; // @[icache.scala 173:46]
  wire  _GEN_441 = io_instAxi_rd_bits_last ? _GEN_312 : _GEN_168; // @[icache.scala 173:46]
  wire  _GEN_442 = io_instAxi_rd_bits_last ? _GEN_313 : _GEN_169; // @[icache.scala 173:46]
  wire  _GEN_443 = io_instAxi_rd_bits_last ? _GEN_314 : _GEN_170; // @[icache.scala 173:46]
  wire  _GEN_444 = io_instAxi_rd_bits_last ? _GEN_315 : _GEN_171; // @[icache.scala 173:46]
  wire  _GEN_445 = io_instAxi_rd_bits_last ? _GEN_316 : _GEN_172; // @[icache.scala 173:46]
  wire  _GEN_446 = io_instAxi_rd_bits_last ? _GEN_317 : _GEN_173; // @[icache.scala 173:46]
  wire  _GEN_447 = io_instAxi_rd_bits_last ? _GEN_318 : _GEN_174; // @[icache.scala 173:46]
  wire  _GEN_448 = io_instAxi_rd_bits_last ? _GEN_319 : _GEN_175; // @[icache.scala 173:46]
  wire  _GEN_449 = io_instAxi_rd_bits_last ? _GEN_320 : _GEN_176; // @[icache.scala 173:46]
  wire  _GEN_450 = io_instAxi_rd_bits_last ? _GEN_321 : _GEN_177; // @[icache.scala 173:46]
  wire  _GEN_451 = io_instAxi_rd_bits_last ? _GEN_322 : _GEN_178; // @[icache.scala 173:46]
  wire  _GEN_452 = io_instAxi_rd_bits_last ? _GEN_323 : _GEN_179; // @[icache.scala 173:46]
  wire  _GEN_453 = io_instAxi_rd_bits_last ? _GEN_324 : _GEN_180; // @[icache.scala 173:46]
  wire  _GEN_454 = io_instAxi_rd_bits_last ? _GEN_325 : _GEN_181; // @[icache.scala 173:46]
  wire  _GEN_455 = io_instAxi_rd_bits_last ? _GEN_326 : _GEN_182; // @[icache.scala 173:46]
  wire  _GEN_456 = io_instAxi_rd_bits_last ? _GEN_327 : _GEN_183; // @[icache.scala 173:46]
  wire  _GEN_457 = io_instAxi_rd_bits_last ? _GEN_328 : _GEN_184; // @[icache.scala 173:46]
  wire  _GEN_458 = io_instAxi_rd_bits_last ? _GEN_329 : _GEN_185; // @[icache.scala 173:46]
  wire  _GEN_459 = io_instAxi_rd_bits_last ? _GEN_330 : _GEN_186; // @[icache.scala 173:46]
  wire  _GEN_460 = io_instAxi_rd_bits_last ? _GEN_331 : _GEN_187; // @[icache.scala 173:46]
  wire  _GEN_461 = io_instAxi_rd_bits_last ? _GEN_332 : _GEN_188; // @[icache.scala 173:46]
  wire  _GEN_462 = io_instAxi_rd_bits_last ? _GEN_333 : _GEN_189; // @[icache.scala 173:46]
  wire  _GEN_463 = io_instAxi_rd_bits_last ? _GEN_334 : _GEN_190; // @[icache.scala 173:46]
  wire  _GEN_464 = io_instAxi_rd_bits_last ? _GEN_335 : _GEN_191; // @[icache.scala 173:46]
  wire  _GEN_465 = io_instAxi_rd_bits_last ? _GEN_336 : _GEN_192; // @[icache.scala 173:46]
  wire  _GEN_466 = io_instAxi_rd_bits_last ? _GEN_337 : _GEN_193; // @[icache.scala 173:46]
  wire [1:0] _GEN_467 = io_instAxi_rd_bits_last ? 2'h0 : state; // @[icache.scala 173:46 icache.scala 177:27 icache.scala 103:24]
  wire [2:0] _GEN_468 = io_instAxi_rd_bits_last ? 3'h0 : _axiOffset_T_1; // @[icache.scala 173:46 icache.scala 178:31 icache.scala 167:27]
  wire [2:0] _GEN_469 = rdataEn & io_instAxi_rd_valid ? _GEN_468 : axiOffset; // @[icache.scala 166:49 icache.scala 81:34]
  wire [63:0] _GEN_471 = rdataEn & io_instAxi_rd_valid ? _GEN_209 : databuf; // @[icache.scala 166:49 icache.scala 82:34]
  wire  _GEN_472 = rdataEn & io_instAxi_rd_valid ? _GEN_338 : rdataEn; // @[icache.scala 166:49 icache.scala 140:30]
  wire [21:0] _GEN_473 = rdataEn & io_instAxi_rd_valid ? _GEN_339 : tag_0_0; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_474 = rdataEn & io_instAxi_rd_valid ? _GEN_340 : tag_0_1; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_475 = rdataEn & io_instAxi_rd_valid ? _GEN_341 : tag_0_2; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_476 = rdataEn & io_instAxi_rd_valid ? _GEN_342 : tag_0_3; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_477 = rdataEn & io_instAxi_rd_valid ? _GEN_343 : tag_0_4; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_478 = rdataEn & io_instAxi_rd_valid ? _GEN_344 : tag_0_5; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_479 = rdataEn & io_instAxi_rd_valid ? _GEN_345 : tag_0_6; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_480 = rdataEn & io_instAxi_rd_valid ? _GEN_346 : tag_0_7; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_481 = rdataEn & io_instAxi_rd_valid ? _GEN_347 : tag_0_8; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_482 = rdataEn & io_instAxi_rd_valid ? _GEN_348 : tag_0_9; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_483 = rdataEn & io_instAxi_rd_valid ? _GEN_349 : tag_0_10; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_484 = rdataEn & io_instAxi_rd_valid ? _GEN_350 : tag_0_11; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_485 = rdataEn & io_instAxi_rd_valid ? _GEN_351 : tag_0_12; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_486 = rdataEn & io_instAxi_rd_valid ? _GEN_352 : tag_0_13; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_487 = rdataEn & io_instAxi_rd_valid ? _GEN_353 : tag_0_14; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_488 = rdataEn & io_instAxi_rd_valid ? _GEN_354 : tag_0_15; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_489 = rdataEn & io_instAxi_rd_valid ? _GEN_355 : tag_1_0; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_490 = rdataEn & io_instAxi_rd_valid ? _GEN_356 : tag_1_1; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_491 = rdataEn & io_instAxi_rd_valid ? _GEN_357 : tag_1_2; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_492 = rdataEn & io_instAxi_rd_valid ? _GEN_358 : tag_1_3; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_493 = rdataEn & io_instAxi_rd_valid ? _GEN_359 : tag_1_4; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_494 = rdataEn & io_instAxi_rd_valid ? _GEN_360 : tag_1_5; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_495 = rdataEn & io_instAxi_rd_valid ? _GEN_361 : tag_1_6; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_496 = rdataEn & io_instAxi_rd_valid ? _GEN_362 : tag_1_7; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_497 = rdataEn & io_instAxi_rd_valid ? _GEN_363 : tag_1_8; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_498 = rdataEn & io_instAxi_rd_valid ? _GEN_364 : tag_1_9; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_499 = rdataEn & io_instAxi_rd_valid ? _GEN_365 : tag_1_10; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_500 = rdataEn & io_instAxi_rd_valid ? _GEN_366 : tag_1_11; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_501 = rdataEn & io_instAxi_rd_valid ? _GEN_367 : tag_1_12; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_502 = rdataEn & io_instAxi_rd_valid ? _GEN_368 : tag_1_13; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_503 = rdataEn & io_instAxi_rd_valid ? _GEN_369 : tag_1_14; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_504 = rdataEn & io_instAxi_rd_valid ? _GEN_370 : tag_1_15; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_505 = rdataEn & io_instAxi_rd_valid ? _GEN_371 : tag_2_0; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_506 = rdataEn & io_instAxi_rd_valid ? _GEN_372 : tag_2_1; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_507 = rdataEn & io_instAxi_rd_valid ? _GEN_373 : tag_2_2; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_508 = rdataEn & io_instAxi_rd_valid ? _GEN_374 : tag_2_3; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_509 = rdataEn & io_instAxi_rd_valid ? _GEN_375 : tag_2_4; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_510 = rdataEn & io_instAxi_rd_valid ? _GEN_376 : tag_2_5; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_511 = rdataEn & io_instAxi_rd_valid ? _GEN_377 : tag_2_6; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_512 = rdataEn & io_instAxi_rd_valid ? _GEN_378 : tag_2_7; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_513 = rdataEn & io_instAxi_rd_valid ? _GEN_379 : tag_2_8; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_514 = rdataEn & io_instAxi_rd_valid ? _GEN_380 : tag_2_9; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_515 = rdataEn & io_instAxi_rd_valid ? _GEN_381 : tag_2_10; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_516 = rdataEn & io_instAxi_rd_valid ? _GEN_382 : tag_2_11; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_517 = rdataEn & io_instAxi_rd_valid ? _GEN_383 : tag_2_12; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_518 = rdataEn & io_instAxi_rd_valid ? _GEN_384 : tag_2_13; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_519 = rdataEn & io_instAxi_rd_valid ? _GEN_385 : tag_2_14; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_520 = rdataEn & io_instAxi_rd_valid ? _GEN_386 : tag_2_15; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_521 = rdataEn & io_instAxi_rd_valid ? _GEN_387 : tag_3_0; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_522 = rdataEn & io_instAxi_rd_valid ? _GEN_388 : tag_3_1; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_523 = rdataEn & io_instAxi_rd_valid ? _GEN_389 : tag_3_2; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_524 = rdataEn & io_instAxi_rd_valid ? _GEN_390 : tag_3_3; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_525 = rdataEn & io_instAxi_rd_valid ? _GEN_391 : tag_3_4; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_526 = rdataEn & io_instAxi_rd_valid ? _GEN_392 : tag_3_5; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_527 = rdataEn & io_instAxi_rd_valid ? _GEN_393 : tag_3_6; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_528 = rdataEn & io_instAxi_rd_valid ? _GEN_394 : tag_3_7; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_529 = rdataEn & io_instAxi_rd_valid ? _GEN_395 : tag_3_8; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_530 = rdataEn & io_instAxi_rd_valid ? _GEN_396 : tag_3_9; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_531 = rdataEn & io_instAxi_rd_valid ? _GEN_397 : tag_3_10; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_532 = rdataEn & io_instAxi_rd_valid ? _GEN_398 : tag_3_11; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_533 = rdataEn & io_instAxi_rd_valid ? _GEN_399 : tag_3_12; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_534 = rdataEn & io_instAxi_rd_valid ? _GEN_400 : tag_3_13; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_535 = rdataEn & io_instAxi_rd_valid ? _GEN_401 : tag_3_14; // @[icache.scala 166:49 icache.scala 69:26]
  wire [21:0] _GEN_536 = rdataEn & io_instAxi_rd_valid ? _GEN_402 : tag_3_15; // @[icache.scala 166:49 icache.scala 69:26]
  wire  _GEN_537 = rdataEn & io_instAxi_rd_valid ? _GEN_403 : _GEN_130; // @[icache.scala 166:49]
  wire  _GEN_538 = rdataEn & io_instAxi_rd_valid ? _GEN_404 : _GEN_131; // @[icache.scala 166:49]
  wire  _GEN_539 = rdataEn & io_instAxi_rd_valid ? _GEN_405 : _GEN_132; // @[icache.scala 166:49]
  wire  _GEN_540 = rdataEn & io_instAxi_rd_valid ? _GEN_406 : _GEN_133; // @[icache.scala 166:49]
  wire  _GEN_541 = rdataEn & io_instAxi_rd_valid ? _GEN_407 : _GEN_134; // @[icache.scala 166:49]
  wire  _GEN_542 = rdataEn & io_instAxi_rd_valid ? _GEN_408 : _GEN_135; // @[icache.scala 166:49]
  wire  _GEN_543 = rdataEn & io_instAxi_rd_valid ? _GEN_409 : _GEN_136; // @[icache.scala 166:49]
  wire  _GEN_544 = rdataEn & io_instAxi_rd_valid ? _GEN_410 : _GEN_137; // @[icache.scala 166:49]
  wire  _GEN_545 = rdataEn & io_instAxi_rd_valid ? _GEN_411 : _GEN_138; // @[icache.scala 166:49]
  wire  _GEN_546 = rdataEn & io_instAxi_rd_valid ? _GEN_412 : _GEN_139; // @[icache.scala 166:49]
  wire  _GEN_547 = rdataEn & io_instAxi_rd_valid ? _GEN_413 : _GEN_140; // @[icache.scala 166:49]
  wire  _GEN_548 = rdataEn & io_instAxi_rd_valid ? _GEN_414 : _GEN_141; // @[icache.scala 166:49]
  wire  _GEN_549 = rdataEn & io_instAxi_rd_valid ? _GEN_415 : _GEN_142; // @[icache.scala 166:49]
  wire  _GEN_550 = rdataEn & io_instAxi_rd_valid ? _GEN_416 : _GEN_143; // @[icache.scala 166:49]
  wire  _GEN_551 = rdataEn & io_instAxi_rd_valid ? _GEN_417 : _GEN_144; // @[icache.scala 166:49]
  wire  _GEN_552 = rdataEn & io_instAxi_rd_valid ? _GEN_418 : _GEN_145; // @[icache.scala 166:49]
  wire  _GEN_553 = rdataEn & io_instAxi_rd_valid ? _GEN_419 : _GEN_146; // @[icache.scala 166:49]
  wire  _GEN_554 = rdataEn & io_instAxi_rd_valid ? _GEN_420 : _GEN_147; // @[icache.scala 166:49]
  wire  _GEN_555 = rdataEn & io_instAxi_rd_valid ? _GEN_421 : _GEN_148; // @[icache.scala 166:49]
  wire  _GEN_556 = rdataEn & io_instAxi_rd_valid ? _GEN_422 : _GEN_149; // @[icache.scala 166:49]
  wire  _GEN_557 = rdataEn & io_instAxi_rd_valid ? _GEN_423 : _GEN_150; // @[icache.scala 166:49]
  wire  _GEN_558 = rdataEn & io_instAxi_rd_valid ? _GEN_424 : _GEN_151; // @[icache.scala 166:49]
  wire  _GEN_559 = rdataEn & io_instAxi_rd_valid ? _GEN_425 : _GEN_152; // @[icache.scala 166:49]
  wire  _GEN_560 = rdataEn & io_instAxi_rd_valid ? _GEN_426 : _GEN_153; // @[icache.scala 166:49]
  wire  _GEN_561 = rdataEn & io_instAxi_rd_valid ? _GEN_427 : _GEN_154; // @[icache.scala 166:49]
  wire  _GEN_562 = rdataEn & io_instAxi_rd_valid ? _GEN_428 : _GEN_155; // @[icache.scala 166:49]
  wire  _GEN_563 = rdataEn & io_instAxi_rd_valid ? _GEN_429 : _GEN_156; // @[icache.scala 166:49]
  wire  _GEN_564 = rdataEn & io_instAxi_rd_valid ? _GEN_430 : _GEN_157; // @[icache.scala 166:49]
  wire  _GEN_565 = rdataEn & io_instAxi_rd_valid ? _GEN_431 : _GEN_158; // @[icache.scala 166:49]
  wire  _GEN_566 = rdataEn & io_instAxi_rd_valid ? _GEN_432 : _GEN_159; // @[icache.scala 166:49]
  wire  _GEN_567 = rdataEn & io_instAxi_rd_valid ? _GEN_433 : _GEN_160; // @[icache.scala 166:49]
  wire  _GEN_568 = rdataEn & io_instAxi_rd_valid ? _GEN_434 : _GEN_161; // @[icache.scala 166:49]
  wire  _GEN_569 = rdataEn & io_instAxi_rd_valid ? _GEN_435 : _GEN_162; // @[icache.scala 166:49]
  wire  _GEN_570 = rdataEn & io_instAxi_rd_valid ? _GEN_436 : _GEN_163; // @[icache.scala 166:49]
  wire  _GEN_571 = rdataEn & io_instAxi_rd_valid ? _GEN_437 : _GEN_164; // @[icache.scala 166:49]
  wire  _GEN_572 = rdataEn & io_instAxi_rd_valid ? _GEN_438 : _GEN_165; // @[icache.scala 166:49]
  wire  _GEN_573 = rdataEn & io_instAxi_rd_valid ? _GEN_439 : _GEN_166; // @[icache.scala 166:49]
  wire  _GEN_574 = rdataEn & io_instAxi_rd_valid ? _GEN_440 : _GEN_167; // @[icache.scala 166:49]
  wire  _GEN_575 = rdataEn & io_instAxi_rd_valid ? _GEN_441 : _GEN_168; // @[icache.scala 166:49]
  wire  _GEN_576 = rdataEn & io_instAxi_rd_valid ? _GEN_442 : _GEN_169; // @[icache.scala 166:49]
  wire  _GEN_577 = rdataEn & io_instAxi_rd_valid ? _GEN_443 : _GEN_170; // @[icache.scala 166:49]
  wire  _GEN_578 = rdataEn & io_instAxi_rd_valid ? _GEN_444 : _GEN_171; // @[icache.scala 166:49]
  wire  _GEN_579 = rdataEn & io_instAxi_rd_valid ? _GEN_445 : _GEN_172; // @[icache.scala 166:49]
  wire  _GEN_580 = rdataEn & io_instAxi_rd_valid ? _GEN_446 : _GEN_173; // @[icache.scala 166:49]
  wire  _GEN_581 = rdataEn & io_instAxi_rd_valid ? _GEN_447 : _GEN_174; // @[icache.scala 166:49]
  wire  _GEN_582 = rdataEn & io_instAxi_rd_valid ? _GEN_448 : _GEN_175; // @[icache.scala 166:49]
  wire  _GEN_583 = rdataEn & io_instAxi_rd_valid ? _GEN_449 : _GEN_176; // @[icache.scala 166:49]
  wire  _GEN_584 = rdataEn & io_instAxi_rd_valid ? _GEN_450 : _GEN_177; // @[icache.scala 166:49]
  wire  _GEN_585 = rdataEn & io_instAxi_rd_valid ? _GEN_451 : _GEN_178; // @[icache.scala 166:49]
  wire  _GEN_586 = rdataEn & io_instAxi_rd_valid ? _GEN_452 : _GEN_179; // @[icache.scala 166:49]
  wire  _GEN_587 = rdataEn & io_instAxi_rd_valid ? _GEN_453 : _GEN_180; // @[icache.scala 166:49]
  wire  _GEN_588 = rdataEn & io_instAxi_rd_valid ? _GEN_454 : _GEN_181; // @[icache.scala 166:49]
  wire  _GEN_589 = rdataEn & io_instAxi_rd_valid ? _GEN_455 : _GEN_182; // @[icache.scala 166:49]
  wire  _GEN_590 = rdataEn & io_instAxi_rd_valid ? _GEN_456 : _GEN_183; // @[icache.scala 166:49]
  wire  _GEN_591 = rdataEn & io_instAxi_rd_valid ? _GEN_457 : _GEN_184; // @[icache.scala 166:49]
  wire  _GEN_592 = rdataEn & io_instAxi_rd_valid ? _GEN_458 : _GEN_185; // @[icache.scala 166:49]
  wire  _GEN_593 = rdataEn & io_instAxi_rd_valid ? _GEN_459 : _GEN_186; // @[icache.scala 166:49]
  wire  _GEN_594 = rdataEn & io_instAxi_rd_valid ? _GEN_460 : _GEN_187; // @[icache.scala 166:49]
  wire  _GEN_595 = rdataEn & io_instAxi_rd_valid ? _GEN_461 : _GEN_188; // @[icache.scala 166:49]
  wire  _GEN_596 = rdataEn & io_instAxi_rd_valid ? _GEN_462 : _GEN_189; // @[icache.scala 166:49]
  wire  _GEN_597 = rdataEn & io_instAxi_rd_valid ? _GEN_463 : _GEN_190; // @[icache.scala 166:49]
  wire  _GEN_598 = rdataEn & io_instAxi_rd_valid ? _GEN_464 : _GEN_191; // @[icache.scala 166:49]
  wire  _GEN_599 = rdataEn & io_instAxi_rd_valid ? _GEN_465 : _GEN_192; // @[icache.scala 166:49]
  wire  _GEN_600 = rdataEn & io_instAxi_rd_valid ? _GEN_466 : _GEN_193; // @[icache.scala 166:49]
  wire [1:0] _GEN_601 = rdataEn & io_instAxi_rd_valid ? _GEN_467 : state; // @[icache.scala 166:49 icache.scala 103:24]
  wire  _GEN_869 = _T & _GEN_199; // @[Conditional.scala 40:58 icache.scala 74:13]
  ysyx_210539_MaxPeriodFibonacciLFSR matchWay_prng ( // @[PRNG.scala 82:22]
    .clock(matchWay_prng_clock),
    .reset(matchWay_prng_reset),
    .io_out_0(matchWay_prng_io_out_0),
    .io_out_1(matchWay_prng_io_out_1),
    .io_out_2(matchWay_prng_io_out_2)
  );
  assign io_instAxi_ra_valid = raddrEn; // @[icache.scala 186:30]
  assign io_instAxi_ra_bits_addr = raddr; // @[icache.scala 187:30]
  assign io_icRead_inst = addr_r[3] ? rdata128[127:64] : rdata128[63:0]; // @[Mux.scala 80:57]
  assign io_icRead_ready = valid_in & ~wait_r; // @[icache.scala 77:37]
  assign io_icRead_rvalid = valid_r; // @[icache.scala 78:25]
  assign io_ic2sr0_addr = state == 2'h2 ? cur_raddr : cur_ram_addr; // @[icache.scala 116:26]
  assign io_ic2sr0_cen = ~(cur_way == 32'h0 & (wait_r | hs_in)); // @[icache.scala 120:23]
  assign io_ic2sr0_wen = ~wen; // @[icache.scala 132:22]
  assign io_ic2sr0_wmask = 128'h0; // @[icache.scala 128:24]
  assign io_ic2sr0_wdata = {io_instAxi_rd_bits_data,databuf}; // @[Cat.scala 30:58]
  assign io_ic2sr1_addr = io_ic2sr0_addr; // @[icache.scala 117:20]
  assign io_ic2sr1_cen = ~(cur_way == 32'h1 & _io_ic2sr0_cen_T_1); // @[icache.scala 121:23]
  assign io_ic2sr1_wen = io_ic2sr0_wen; // @[icache.scala 133:19]
  assign io_ic2sr1_wmask = io_ic2sr0_wmask; // @[icache.scala 129:21]
  assign io_ic2sr1_wdata = io_ic2sr0_wdata; // @[icache.scala 125:21]
  assign io_ic2sr2_addr = io_ic2sr0_addr; // @[icache.scala 118:20]
  assign io_ic2sr2_cen = ~(cur_way == 32'h2 & _io_ic2sr0_cen_T_1); // @[icache.scala 122:23]
  assign io_ic2sr2_wen = io_ic2sr0_wen; // @[icache.scala 134:19]
  assign io_ic2sr2_wmask = io_ic2sr0_wmask; // @[icache.scala 130:21]
  assign io_ic2sr2_wdata = io_ic2sr0_wdata; // @[icache.scala 126:21]
  assign io_ic2sr3_addr = io_ic2sr0_addr; // @[icache.scala 119:20]
  assign io_ic2sr3_cen = ~(cur_way == 32'h3 & _io_ic2sr0_cen_T_1); // @[icache.scala 123:23]
  assign io_ic2sr3_wen = io_ic2sr0_wen; // @[icache.scala 135:19]
  assign io_ic2sr3_wmask = io_ic2sr0_wmask; // @[icache.scala 131:21]
  assign io_ic2sr3_wdata = io_ic2sr0_wdata; // @[icache.scala 127:21]
  assign matchWay_prng_clock = clock;
  assign matchWay_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[icache.scala 69:26]
      tag_0_0 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_0_0 <= _GEN_473;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_0_1 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_0_1 <= _GEN_474;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_0_2 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_0_2 <= _GEN_475;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_0_3 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_0_3 <= _GEN_476;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_0_4 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_0_4 <= _GEN_477;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_0_5 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_0_5 <= _GEN_478;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_0_6 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_0_6 <= _GEN_479;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_0_7 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_0_7 <= _GEN_480;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_0_8 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_0_8 <= _GEN_481;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_0_9 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_0_9 <= _GEN_482;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_0_10 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_0_10 <= _GEN_483;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_0_11 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_0_11 <= _GEN_484;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_0_12 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_0_12 <= _GEN_485;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_0_13 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_0_13 <= _GEN_486;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_0_14 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_0_14 <= _GEN_487;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_0_15 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_0_15 <= _GEN_488;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_1_0 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_1_0 <= _GEN_489;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_1_1 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_1_1 <= _GEN_490;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_1_2 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_1_2 <= _GEN_491;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_1_3 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_1_3 <= _GEN_492;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_1_4 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_1_4 <= _GEN_493;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_1_5 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_1_5 <= _GEN_494;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_1_6 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_1_6 <= _GEN_495;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_1_7 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_1_7 <= _GEN_496;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_1_8 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_1_8 <= _GEN_497;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_1_9 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_1_9 <= _GEN_498;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_1_10 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_1_10 <= _GEN_499;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_1_11 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_1_11 <= _GEN_500;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_1_12 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_1_12 <= _GEN_501;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_1_13 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_1_13 <= _GEN_502;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_1_14 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_1_14 <= _GEN_503;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_1_15 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_1_15 <= _GEN_504;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_2_0 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_2_0 <= _GEN_505;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_2_1 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_2_1 <= _GEN_506;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_2_2 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_2_2 <= _GEN_507;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_2_3 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_2_3 <= _GEN_508;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_2_4 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_2_4 <= _GEN_509;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_2_5 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_2_5 <= _GEN_510;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_2_6 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_2_6 <= _GEN_511;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_2_7 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_2_7 <= _GEN_512;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_2_8 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_2_8 <= _GEN_513;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_2_9 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_2_9 <= _GEN_514;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_2_10 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_2_10 <= _GEN_515;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_2_11 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_2_11 <= _GEN_516;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_2_12 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_2_12 <= _GEN_517;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_2_13 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_2_13 <= _GEN_518;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_2_14 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_2_14 <= _GEN_519;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_2_15 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_2_15 <= _GEN_520;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_3_0 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_3_0 <= _GEN_521;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_3_1 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_3_1 <= _GEN_522;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_3_2 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_3_2 <= _GEN_523;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_3_3 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_3_3 <= _GEN_524;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_3_4 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_3_4 <= _GEN_525;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_3_5 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_3_5 <= _GEN_526;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_3_6 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_3_6 <= _GEN_527;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_3_7 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_3_7 <= _GEN_528;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_3_8 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_3_8 <= _GEN_529;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_3_9 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_3_9 <= _GEN_530;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_3_10 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_3_10 <= _GEN_531;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_3_11 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_3_11 <= _GEN_532;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_3_12 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_3_12 <= _GEN_533;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_3_13 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_3_13 <= _GEN_534;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_3_14 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_3_14 <= _GEN_535;
        end
      end
    end
    if (reset) begin // @[icache.scala 69:26]
      tag_3_15 <= 22'h0; // @[icache.scala 69:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          tag_3_15 <= _GEN_536;
        end
      end
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_0_0 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_0_0 <= _GEN_130;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_0_0 <= _GEN_130;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_0_0 <= _GEN_537;
    end else begin
      valid_0_0 <= _GEN_130;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_0_1 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_0_1 <= _GEN_131;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_0_1 <= _GEN_131;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_0_1 <= _GEN_538;
    end else begin
      valid_0_1 <= _GEN_131;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_0_2 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_0_2 <= _GEN_132;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_0_2 <= _GEN_132;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_0_2 <= _GEN_539;
    end else begin
      valid_0_2 <= _GEN_132;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_0_3 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_0_3 <= _GEN_133;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_0_3 <= _GEN_133;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_0_3 <= _GEN_540;
    end else begin
      valid_0_3 <= _GEN_133;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_0_4 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_0_4 <= _GEN_134;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_0_4 <= _GEN_134;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_0_4 <= _GEN_541;
    end else begin
      valid_0_4 <= _GEN_134;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_0_5 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_0_5 <= _GEN_135;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_0_5 <= _GEN_135;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_0_5 <= _GEN_542;
    end else begin
      valid_0_5 <= _GEN_135;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_0_6 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_0_6 <= _GEN_136;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_0_6 <= _GEN_136;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_0_6 <= _GEN_543;
    end else begin
      valid_0_6 <= _GEN_136;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_0_7 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_0_7 <= _GEN_137;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_0_7 <= _GEN_137;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_0_7 <= _GEN_544;
    end else begin
      valid_0_7 <= _GEN_137;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_0_8 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_0_8 <= _GEN_138;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_0_8 <= _GEN_138;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_0_8 <= _GEN_545;
    end else begin
      valid_0_8 <= _GEN_138;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_0_9 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_0_9 <= _GEN_139;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_0_9 <= _GEN_139;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_0_9 <= _GEN_546;
    end else begin
      valid_0_9 <= _GEN_139;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_0_10 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_0_10 <= _GEN_140;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_0_10 <= _GEN_140;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_0_10 <= _GEN_547;
    end else begin
      valid_0_10 <= _GEN_140;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_0_11 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_0_11 <= _GEN_141;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_0_11 <= _GEN_141;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_0_11 <= _GEN_548;
    end else begin
      valid_0_11 <= _GEN_141;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_0_12 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_0_12 <= _GEN_142;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_0_12 <= _GEN_142;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_0_12 <= _GEN_549;
    end else begin
      valid_0_12 <= _GEN_142;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_0_13 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_0_13 <= _GEN_143;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_0_13 <= _GEN_143;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_0_13 <= _GEN_550;
    end else begin
      valid_0_13 <= _GEN_143;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_0_14 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_0_14 <= _GEN_144;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_0_14 <= _GEN_144;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_0_14 <= _GEN_551;
    end else begin
      valid_0_14 <= _GEN_144;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_0_15 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_0_15 <= _GEN_145;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_0_15 <= _GEN_145;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_0_15 <= _GEN_552;
    end else begin
      valid_0_15 <= _GEN_145;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_1_0 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_1_0 <= _GEN_146;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_1_0 <= _GEN_146;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_1_0 <= _GEN_553;
    end else begin
      valid_1_0 <= _GEN_146;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_1_1 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_1_1 <= _GEN_147;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_1_1 <= _GEN_147;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_1_1 <= _GEN_554;
    end else begin
      valid_1_1 <= _GEN_147;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_1_2 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_1_2 <= _GEN_148;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_1_2 <= _GEN_148;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_1_2 <= _GEN_555;
    end else begin
      valid_1_2 <= _GEN_148;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_1_3 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_1_3 <= _GEN_149;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_1_3 <= _GEN_149;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_1_3 <= _GEN_556;
    end else begin
      valid_1_3 <= _GEN_149;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_1_4 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_1_4 <= _GEN_150;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_1_4 <= _GEN_150;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_1_4 <= _GEN_557;
    end else begin
      valid_1_4 <= _GEN_150;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_1_5 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_1_5 <= _GEN_151;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_1_5 <= _GEN_151;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_1_5 <= _GEN_558;
    end else begin
      valid_1_5 <= _GEN_151;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_1_6 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_1_6 <= _GEN_152;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_1_6 <= _GEN_152;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_1_6 <= _GEN_559;
    end else begin
      valid_1_6 <= _GEN_152;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_1_7 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_1_7 <= _GEN_153;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_1_7 <= _GEN_153;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_1_7 <= _GEN_560;
    end else begin
      valid_1_7 <= _GEN_153;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_1_8 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_1_8 <= _GEN_154;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_1_8 <= _GEN_154;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_1_8 <= _GEN_561;
    end else begin
      valid_1_8 <= _GEN_154;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_1_9 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_1_9 <= _GEN_155;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_1_9 <= _GEN_155;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_1_9 <= _GEN_562;
    end else begin
      valid_1_9 <= _GEN_155;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_1_10 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_1_10 <= _GEN_156;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_1_10 <= _GEN_156;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_1_10 <= _GEN_563;
    end else begin
      valid_1_10 <= _GEN_156;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_1_11 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_1_11 <= _GEN_157;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_1_11 <= _GEN_157;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_1_11 <= _GEN_564;
    end else begin
      valid_1_11 <= _GEN_157;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_1_12 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_1_12 <= _GEN_158;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_1_12 <= _GEN_158;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_1_12 <= _GEN_565;
    end else begin
      valid_1_12 <= _GEN_158;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_1_13 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_1_13 <= _GEN_159;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_1_13 <= _GEN_159;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_1_13 <= _GEN_566;
    end else begin
      valid_1_13 <= _GEN_159;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_1_14 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_1_14 <= _GEN_160;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_1_14 <= _GEN_160;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_1_14 <= _GEN_567;
    end else begin
      valid_1_14 <= _GEN_160;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_1_15 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_1_15 <= _GEN_161;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_1_15 <= _GEN_161;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_1_15 <= _GEN_568;
    end else begin
      valid_1_15 <= _GEN_161;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_2_0 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_2_0 <= _GEN_162;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_2_0 <= _GEN_162;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_2_0 <= _GEN_569;
    end else begin
      valid_2_0 <= _GEN_162;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_2_1 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_2_1 <= _GEN_163;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_2_1 <= _GEN_163;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_2_1 <= _GEN_570;
    end else begin
      valid_2_1 <= _GEN_163;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_2_2 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_2_2 <= _GEN_164;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_2_2 <= _GEN_164;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_2_2 <= _GEN_571;
    end else begin
      valid_2_2 <= _GEN_164;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_2_3 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_2_3 <= _GEN_165;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_2_3 <= _GEN_165;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_2_3 <= _GEN_572;
    end else begin
      valid_2_3 <= _GEN_165;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_2_4 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_2_4 <= _GEN_166;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_2_4 <= _GEN_166;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_2_4 <= _GEN_573;
    end else begin
      valid_2_4 <= _GEN_166;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_2_5 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_2_5 <= _GEN_167;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_2_5 <= _GEN_167;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_2_5 <= _GEN_574;
    end else begin
      valid_2_5 <= _GEN_167;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_2_6 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_2_6 <= _GEN_168;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_2_6 <= _GEN_168;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_2_6 <= _GEN_575;
    end else begin
      valid_2_6 <= _GEN_168;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_2_7 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_2_7 <= _GEN_169;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_2_7 <= _GEN_169;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_2_7 <= _GEN_576;
    end else begin
      valid_2_7 <= _GEN_169;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_2_8 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_2_8 <= _GEN_170;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_2_8 <= _GEN_170;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_2_8 <= _GEN_577;
    end else begin
      valid_2_8 <= _GEN_170;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_2_9 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_2_9 <= _GEN_171;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_2_9 <= _GEN_171;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_2_9 <= _GEN_578;
    end else begin
      valid_2_9 <= _GEN_171;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_2_10 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_2_10 <= _GEN_172;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_2_10 <= _GEN_172;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_2_10 <= _GEN_579;
    end else begin
      valid_2_10 <= _GEN_172;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_2_11 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_2_11 <= _GEN_173;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_2_11 <= _GEN_173;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_2_11 <= _GEN_580;
    end else begin
      valid_2_11 <= _GEN_173;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_2_12 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_2_12 <= _GEN_174;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_2_12 <= _GEN_174;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_2_12 <= _GEN_581;
    end else begin
      valid_2_12 <= _GEN_174;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_2_13 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_2_13 <= _GEN_175;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_2_13 <= _GEN_175;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_2_13 <= _GEN_582;
    end else begin
      valid_2_13 <= _GEN_175;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_2_14 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_2_14 <= _GEN_176;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_2_14 <= _GEN_176;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_2_14 <= _GEN_583;
    end else begin
      valid_2_14 <= _GEN_176;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_2_15 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_2_15 <= _GEN_177;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_2_15 <= _GEN_177;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_2_15 <= _GEN_584;
    end else begin
      valid_2_15 <= _GEN_177;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_3_0 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_3_0 <= _GEN_178;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_3_0 <= _GEN_178;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_3_0 <= _GEN_585;
    end else begin
      valid_3_0 <= _GEN_178;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_3_1 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_3_1 <= _GEN_179;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_3_1 <= _GEN_179;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_3_1 <= _GEN_586;
    end else begin
      valid_3_1 <= _GEN_179;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_3_2 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_3_2 <= _GEN_180;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_3_2 <= _GEN_180;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_3_2 <= _GEN_587;
    end else begin
      valid_3_2 <= _GEN_180;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_3_3 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_3_3 <= _GEN_181;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_3_3 <= _GEN_181;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_3_3 <= _GEN_588;
    end else begin
      valid_3_3 <= _GEN_181;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_3_4 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_3_4 <= _GEN_182;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_3_4 <= _GEN_182;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_3_4 <= _GEN_589;
    end else begin
      valid_3_4 <= _GEN_182;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_3_5 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_3_5 <= _GEN_183;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_3_5 <= _GEN_183;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_3_5 <= _GEN_590;
    end else begin
      valid_3_5 <= _GEN_183;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_3_6 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_3_6 <= _GEN_184;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_3_6 <= _GEN_184;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_3_6 <= _GEN_591;
    end else begin
      valid_3_6 <= _GEN_184;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_3_7 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_3_7 <= _GEN_185;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_3_7 <= _GEN_185;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_3_7 <= _GEN_592;
    end else begin
      valid_3_7 <= _GEN_185;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_3_8 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_3_8 <= _GEN_186;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_3_8 <= _GEN_186;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_3_8 <= _GEN_593;
    end else begin
      valid_3_8 <= _GEN_186;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_3_9 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_3_9 <= _GEN_187;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_3_9 <= _GEN_187;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_3_9 <= _GEN_594;
    end else begin
      valid_3_9 <= _GEN_187;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_3_10 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_3_10 <= _GEN_188;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_3_10 <= _GEN_188;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_3_10 <= _GEN_595;
    end else begin
      valid_3_10 <= _GEN_188;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_3_11 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_3_11 <= _GEN_189;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_3_11 <= _GEN_189;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_3_11 <= _GEN_596;
    end else begin
      valid_3_11 <= _GEN_189;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_3_12 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_3_12 <= _GEN_190;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_3_12 <= _GEN_190;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_3_12 <= _GEN_597;
    end else begin
      valid_3_12 <= _GEN_190;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_3_13 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_3_13 <= _GEN_191;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_3_13 <= _GEN_191;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_3_13 <= _GEN_598;
    end else begin
      valid_3_13 <= _GEN_191;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_3_14 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_3_14 <= _GEN_192;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_3_14 <= _GEN_192;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_3_14 <= _GEN_599;
    end else begin
      valid_3_14 <= _GEN_192;
    end
    if (reset) begin // @[icache.scala 70:26]
      valid_3_15 <= 1'h0; // @[icache.scala 70:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      valid_3_15 <= _GEN_193;
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      valid_3_15 <= _GEN_193;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      valid_3_15 <= _GEN_600;
    end else begin
      valid_3_15 <= _GEN_193;
    end
    if (reset) begin // @[icache.scala 72:30]
      wait_r <= 1'h0; // @[icache.scala 72:30]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (!(~hs_in & _io_icRead_ready_T)) begin // @[icache.scala 144:36]
        if (cacheHit) begin // @[icache.scala 146:33]
          wait_r <= 1'h0; // @[icache.scala 148:25]
        end else begin
          wait_r <= 1'h1; // @[icache.scala 154:25]
        end
      end
    end
    if (reset) begin // @[icache.scala 73:30]
      valid_r <= 1'h0; // @[icache.scala 73:30]
    end else begin
      valid_r <= _GEN_869;
    end
    if (reset) begin // @[icache.scala 79:34]
      addr_r <= 32'h0; // @[icache.scala 79:34]
    end else if (hs_in) begin // @[icache.scala 83:30]
      addr_r <= io_icRead_addr;
    end
    if (reset) begin // @[icache.scala 80:34]
      matchWay_r <= 32'h0; // @[icache.scala 80:34]
    end else if (hs_in) begin // @[icache.scala 91:30]
      matchWay_r <= {{30'd0}, matchWay};
    end
    if (reset) begin // @[icache.scala 81:34]
      axiOffset <= 3'h0; // @[icache.scala 81:34]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_4) begin // @[Conditional.scala 39:67]
        if (raddrEn & io_instAxi_ra_ready) begin // @[icache.scala 158:49]
          axiOffset <= 3'h0; // @[icache.scala 162:27]
        end
      end else if (_T_6) begin // @[Conditional.scala 39:67]
        axiOffset <= _GEN_469;
      end
    end
    if (reset) begin // @[icache.scala 82:34]
      databuf <= 64'h0; // @[icache.scala 82:34]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_4)) begin // @[Conditional.scala 39:67]
        if (_T_6) begin // @[Conditional.scala 39:67]
          databuf <= _GEN_471;
        end
      end
    end
    if (reset) begin // @[icache.scala 103:24]
      state <= 2'h0; // @[icache.scala 103:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (!(~hs_in & _io_icRead_ready_T)) begin // @[icache.scala 144:36]
        if (!(cacheHit)) begin // @[icache.scala 146:33]
          state <= 2'h1; // @[icache.scala 152:25]
        end
      end
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      if (raddrEn & io_instAxi_ra_ready) begin // @[icache.scala 158:49]
        state <= 2'h2; // @[icache.scala 159:25]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      state <= _GEN_601;
    end
    if (reset) begin // @[icache.scala 140:30]
      rdataEn <= 1'h0; // @[icache.scala 140:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_4) begin // @[Conditional.scala 39:67]
        rdataEn <= _GEN_206;
      end else if (_T_6) begin // @[Conditional.scala 39:67]
        rdataEn <= _GEN_472;
      end
    end
    if (reset) begin // @[icache.scala 138:30]
      raddrEn <= 1'h0; // @[icache.scala 138:30]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (!(~hs_in & _io_icRead_ready_T)) begin // @[icache.scala 144:36]
        if (!(cacheHit)) begin // @[icache.scala 146:33]
          raddrEn <= 1'h1; // @[icache.scala 151:25]
        end
      end
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      if (raddrEn & io_instAxi_ra_ready) begin // @[icache.scala 158:49]
        raddrEn <= 1'h0; // @[icache.scala 160:25]
      end
    end
    if (reset) begin // @[icache.scala 139:30]
      raddr <= 32'h0; // @[icache.scala 139:30]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (!(~hs_in & _io_icRead_ready_T)) begin // @[icache.scala 144:36]
        if (!(cacheHit)) begin // @[icache.scala 146:33]
          raddr <= _raddr_T; // @[icache.scala 150:25]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_0_0 = _RAND_0[21:0];
  _RAND_1 = {1{`RANDOM}};
  tag_0_1 = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  tag_0_2 = _RAND_2[21:0];
  _RAND_3 = {1{`RANDOM}};
  tag_0_3 = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  tag_0_4 = _RAND_4[21:0];
  _RAND_5 = {1{`RANDOM}};
  tag_0_5 = _RAND_5[21:0];
  _RAND_6 = {1{`RANDOM}};
  tag_0_6 = _RAND_6[21:0];
  _RAND_7 = {1{`RANDOM}};
  tag_0_7 = _RAND_7[21:0];
  _RAND_8 = {1{`RANDOM}};
  tag_0_8 = _RAND_8[21:0];
  _RAND_9 = {1{`RANDOM}};
  tag_0_9 = _RAND_9[21:0];
  _RAND_10 = {1{`RANDOM}};
  tag_0_10 = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  tag_0_11 = _RAND_11[21:0];
  _RAND_12 = {1{`RANDOM}};
  tag_0_12 = _RAND_12[21:0];
  _RAND_13 = {1{`RANDOM}};
  tag_0_13 = _RAND_13[21:0];
  _RAND_14 = {1{`RANDOM}};
  tag_0_14 = _RAND_14[21:0];
  _RAND_15 = {1{`RANDOM}};
  tag_0_15 = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  tag_1_0 = _RAND_16[21:0];
  _RAND_17 = {1{`RANDOM}};
  tag_1_1 = _RAND_17[21:0];
  _RAND_18 = {1{`RANDOM}};
  tag_1_2 = _RAND_18[21:0];
  _RAND_19 = {1{`RANDOM}};
  tag_1_3 = _RAND_19[21:0];
  _RAND_20 = {1{`RANDOM}};
  tag_1_4 = _RAND_20[21:0];
  _RAND_21 = {1{`RANDOM}};
  tag_1_5 = _RAND_21[21:0];
  _RAND_22 = {1{`RANDOM}};
  tag_1_6 = _RAND_22[21:0];
  _RAND_23 = {1{`RANDOM}};
  tag_1_7 = _RAND_23[21:0];
  _RAND_24 = {1{`RANDOM}};
  tag_1_8 = _RAND_24[21:0];
  _RAND_25 = {1{`RANDOM}};
  tag_1_9 = _RAND_25[21:0];
  _RAND_26 = {1{`RANDOM}};
  tag_1_10 = _RAND_26[21:0];
  _RAND_27 = {1{`RANDOM}};
  tag_1_11 = _RAND_27[21:0];
  _RAND_28 = {1{`RANDOM}};
  tag_1_12 = _RAND_28[21:0];
  _RAND_29 = {1{`RANDOM}};
  tag_1_13 = _RAND_29[21:0];
  _RAND_30 = {1{`RANDOM}};
  tag_1_14 = _RAND_30[21:0];
  _RAND_31 = {1{`RANDOM}};
  tag_1_15 = _RAND_31[21:0];
  _RAND_32 = {1{`RANDOM}};
  tag_2_0 = _RAND_32[21:0];
  _RAND_33 = {1{`RANDOM}};
  tag_2_1 = _RAND_33[21:0];
  _RAND_34 = {1{`RANDOM}};
  tag_2_2 = _RAND_34[21:0];
  _RAND_35 = {1{`RANDOM}};
  tag_2_3 = _RAND_35[21:0];
  _RAND_36 = {1{`RANDOM}};
  tag_2_4 = _RAND_36[21:0];
  _RAND_37 = {1{`RANDOM}};
  tag_2_5 = _RAND_37[21:0];
  _RAND_38 = {1{`RANDOM}};
  tag_2_6 = _RAND_38[21:0];
  _RAND_39 = {1{`RANDOM}};
  tag_2_7 = _RAND_39[21:0];
  _RAND_40 = {1{`RANDOM}};
  tag_2_8 = _RAND_40[21:0];
  _RAND_41 = {1{`RANDOM}};
  tag_2_9 = _RAND_41[21:0];
  _RAND_42 = {1{`RANDOM}};
  tag_2_10 = _RAND_42[21:0];
  _RAND_43 = {1{`RANDOM}};
  tag_2_11 = _RAND_43[21:0];
  _RAND_44 = {1{`RANDOM}};
  tag_2_12 = _RAND_44[21:0];
  _RAND_45 = {1{`RANDOM}};
  tag_2_13 = _RAND_45[21:0];
  _RAND_46 = {1{`RANDOM}};
  tag_2_14 = _RAND_46[21:0];
  _RAND_47 = {1{`RANDOM}};
  tag_2_15 = _RAND_47[21:0];
  _RAND_48 = {1{`RANDOM}};
  tag_3_0 = _RAND_48[21:0];
  _RAND_49 = {1{`RANDOM}};
  tag_3_1 = _RAND_49[21:0];
  _RAND_50 = {1{`RANDOM}};
  tag_3_2 = _RAND_50[21:0];
  _RAND_51 = {1{`RANDOM}};
  tag_3_3 = _RAND_51[21:0];
  _RAND_52 = {1{`RANDOM}};
  tag_3_4 = _RAND_52[21:0];
  _RAND_53 = {1{`RANDOM}};
  tag_3_5 = _RAND_53[21:0];
  _RAND_54 = {1{`RANDOM}};
  tag_3_6 = _RAND_54[21:0];
  _RAND_55 = {1{`RANDOM}};
  tag_3_7 = _RAND_55[21:0];
  _RAND_56 = {1{`RANDOM}};
  tag_3_8 = _RAND_56[21:0];
  _RAND_57 = {1{`RANDOM}};
  tag_3_9 = _RAND_57[21:0];
  _RAND_58 = {1{`RANDOM}};
  tag_3_10 = _RAND_58[21:0];
  _RAND_59 = {1{`RANDOM}};
  tag_3_11 = _RAND_59[21:0];
  _RAND_60 = {1{`RANDOM}};
  tag_3_12 = _RAND_60[21:0];
  _RAND_61 = {1{`RANDOM}};
  tag_3_13 = _RAND_61[21:0];
  _RAND_62 = {1{`RANDOM}};
  tag_3_14 = _RAND_62[21:0];
  _RAND_63 = {1{`RANDOM}};
  tag_3_15 = _RAND_63[21:0];
  _RAND_64 = {1{`RANDOM}};
  valid_0_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_0_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_0_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  valid_0_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  valid_0_4 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  valid_0_5 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  valid_0_6 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  valid_0_7 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  valid_0_8 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  valid_0_9 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  valid_0_10 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid_0_11 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  valid_0_12 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  valid_0_13 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  valid_0_14 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  valid_0_15 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  valid_1_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_1_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_1_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_1_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_1_4 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_1_5 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_1_6 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_1_7 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_1_8 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_1_9 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_1_10 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_1_11 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_1_12 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_1_13 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_1_14 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_1_15 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  valid_2_0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  valid_2_1 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  valid_2_2 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  valid_2_3 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  valid_2_4 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  valid_2_5 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  valid_2_6 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  valid_2_7 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  valid_2_8 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  valid_2_9 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  valid_2_10 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  valid_2_11 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  valid_2_12 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  valid_2_13 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  valid_2_14 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  valid_2_15 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  valid_3_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  valid_3_1 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  valid_3_2 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  valid_3_3 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  valid_3_4 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  valid_3_5 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  valid_3_6 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  valid_3_7 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  valid_3_8 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  valid_3_9 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  valid_3_10 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  valid_3_11 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  valid_3_12 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  valid_3_13 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  valid_3_14 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  valid_3_15 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  wait_r = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_r = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  addr_r = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  matchWay_r = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  axiOffset = _RAND_132[2:0];
  _RAND_133 = {2{`RANDOM}};
  databuf = _RAND_133[63:0];
  _RAND_134 = {1{`RANDOM}};
  state = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  rdataEn = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  raddrEn = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  raddr = _RAND_137[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_DataCache(
  input          clock,
  input          reset,
  input          io_dataAxi_wa_ready,
  output         io_dataAxi_wa_valid,
  output [31:0]  io_dataAxi_wa_bits_addr,
  input          io_dataAxi_wd_ready,
  output         io_dataAxi_wd_valid,
  output [63:0]  io_dataAxi_wd_bits_data,
  output         io_dataAxi_wd_bits_last,
  input          io_dataAxi_ra_ready,
  output         io_dataAxi_ra_valid,
  output [31:0]  io_dataAxi_ra_bits_addr,
  input          io_dataAxi_rd_valid,
  input  [63:0]  io_dataAxi_rd_bits_data,
  input          io_dataAxi_rd_bits_last,
  input  [31:0]  io_dcRW_addr,
  output [63:0]  io_dcRW_rdata,
  output         io_dcRW_rvalid,
  input  [63:0]  io_dcRW_wdata,
  input  [4:0]   io_dcRW_dc_mode,
  input  [4:0]   io_dcRW_amo,
  output         io_dcRW_ready,
  input          io_flush,
  output         io_flush_out,
  output [5:0]   io_dc2sr0_addr,
  output         io_dc2sr0_cen,
  output         io_dc2sr0_wen,
  output [127:0] io_dc2sr0_wmask,
  output [127:0] io_dc2sr0_wdata,
  input  [127:0] io_dc2sr0_rdata,
  output [5:0]   io_dc2sr1_addr,
  output         io_dc2sr1_cen,
  output         io_dc2sr1_wen,
  output [127:0] io_dc2sr1_wmask,
  output [127:0] io_dc2sr1_wdata,
  input  [127:0] io_dc2sr1_rdata,
  output [5:0]   io_dc2sr2_addr,
  output         io_dc2sr2_cen,
  output         io_dc2sr2_wen,
  output [127:0] io_dc2sr2_wmask,
  output [127:0] io_dc2sr2_wdata,
  input  [127:0] io_dc2sr2_rdata,
  output [5:0]   io_dc2sr3_addr,
  output         io_dc2sr3_cen,
  output         io_dc2sr3_wen,
  output [127:0] io_dc2sr3_wmask,
  output [127:0] io_dc2sr3_wdata,
  input  [127:0] io_dc2sr3_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
`endif // RANDOMIZE_REG_INIT
  wire  matchWay_prng_clock; // @[PRNG.scala 82:22]
  wire  matchWay_prng_reset; // @[PRNG.scala 82:22]
  wire  matchWay_prng_io_out_0; // @[PRNG.scala 82:22]
  wire  matchWay_prng_io_out_1; // @[PRNG.scala 82:22]
  wire  matchWay_prng_io_out_2; // @[PRNG.scala 82:22]
  reg [21:0] tag_0_0; // @[dcache.scala 92:26]
  reg [21:0] tag_0_1; // @[dcache.scala 92:26]
  reg [21:0] tag_0_2; // @[dcache.scala 92:26]
  reg [21:0] tag_0_3; // @[dcache.scala 92:26]
  reg [21:0] tag_0_4; // @[dcache.scala 92:26]
  reg [21:0] tag_0_5; // @[dcache.scala 92:26]
  reg [21:0] tag_0_6; // @[dcache.scala 92:26]
  reg [21:0] tag_0_7; // @[dcache.scala 92:26]
  reg [21:0] tag_0_8; // @[dcache.scala 92:26]
  reg [21:0] tag_0_9; // @[dcache.scala 92:26]
  reg [21:0] tag_0_10; // @[dcache.scala 92:26]
  reg [21:0] tag_0_11; // @[dcache.scala 92:26]
  reg [21:0] tag_0_12; // @[dcache.scala 92:26]
  reg [21:0] tag_0_13; // @[dcache.scala 92:26]
  reg [21:0] tag_0_14; // @[dcache.scala 92:26]
  reg [21:0] tag_0_15; // @[dcache.scala 92:26]
  reg [21:0] tag_1_0; // @[dcache.scala 92:26]
  reg [21:0] tag_1_1; // @[dcache.scala 92:26]
  reg [21:0] tag_1_2; // @[dcache.scala 92:26]
  reg [21:0] tag_1_3; // @[dcache.scala 92:26]
  reg [21:0] tag_1_4; // @[dcache.scala 92:26]
  reg [21:0] tag_1_5; // @[dcache.scala 92:26]
  reg [21:0] tag_1_6; // @[dcache.scala 92:26]
  reg [21:0] tag_1_7; // @[dcache.scala 92:26]
  reg [21:0] tag_1_8; // @[dcache.scala 92:26]
  reg [21:0] tag_1_9; // @[dcache.scala 92:26]
  reg [21:0] tag_1_10; // @[dcache.scala 92:26]
  reg [21:0] tag_1_11; // @[dcache.scala 92:26]
  reg [21:0] tag_1_12; // @[dcache.scala 92:26]
  reg [21:0] tag_1_13; // @[dcache.scala 92:26]
  reg [21:0] tag_1_14; // @[dcache.scala 92:26]
  reg [21:0] tag_1_15; // @[dcache.scala 92:26]
  reg [21:0] tag_2_0; // @[dcache.scala 92:26]
  reg [21:0] tag_2_1; // @[dcache.scala 92:26]
  reg [21:0] tag_2_2; // @[dcache.scala 92:26]
  reg [21:0] tag_2_3; // @[dcache.scala 92:26]
  reg [21:0] tag_2_4; // @[dcache.scala 92:26]
  reg [21:0] tag_2_5; // @[dcache.scala 92:26]
  reg [21:0] tag_2_6; // @[dcache.scala 92:26]
  reg [21:0] tag_2_7; // @[dcache.scala 92:26]
  reg [21:0] tag_2_8; // @[dcache.scala 92:26]
  reg [21:0] tag_2_9; // @[dcache.scala 92:26]
  reg [21:0] tag_2_10; // @[dcache.scala 92:26]
  reg [21:0] tag_2_11; // @[dcache.scala 92:26]
  reg [21:0] tag_2_12; // @[dcache.scala 92:26]
  reg [21:0] tag_2_13; // @[dcache.scala 92:26]
  reg [21:0] tag_2_14; // @[dcache.scala 92:26]
  reg [21:0] tag_2_15; // @[dcache.scala 92:26]
  reg [21:0] tag_3_0; // @[dcache.scala 92:26]
  reg [21:0] tag_3_1; // @[dcache.scala 92:26]
  reg [21:0] tag_3_2; // @[dcache.scala 92:26]
  reg [21:0] tag_3_3; // @[dcache.scala 92:26]
  reg [21:0] tag_3_4; // @[dcache.scala 92:26]
  reg [21:0] tag_3_5; // @[dcache.scala 92:26]
  reg [21:0] tag_3_6; // @[dcache.scala 92:26]
  reg [21:0] tag_3_7; // @[dcache.scala 92:26]
  reg [21:0] tag_3_8; // @[dcache.scala 92:26]
  reg [21:0] tag_3_9; // @[dcache.scala 92:26]
  reg [21:0] tag_3_10; // @[dcache.scala 92:26]
  reg [21:0] tag_3_11; // @[dcache.scala 92:26]
  reg [21:0] tag_3_12; // @[dcache.scala 92:26]
  reg [21:0] tag_3_13; // @[dcache.scala 92:26]
  reg [21:0] tag_3_14; // @[dcache.scala 92:26]
  reg [21:0] tag_3_15; // @[dcache.scala 92:26]
  reg  valid_0_0; // @[dcache.scala 93:26]
  reg  valid_0_1; // @[dcache.scala 93:26]
  reg  valid_0_2; // @[dcache.scala 93:26]
  reg  valid_0_3; // @[dcache.scala 93:26]
  reg  valid_0_4; // @[dcache.scala 93:26]
  reg  valid_0_5; // @[dcache.scala 93:26]
  reg  valid_0_6; // @[dcache.scala 93:26]
  reg  valid_0_7; // @[dcache.scala 93:26]
  reg  valid_0_8; // @[dcache.scala 93:26]
  reg  valid_0_9; // @[dcache.scala 93:26]
  reg  valid_0_10; // @[dcache.scala 93:26]
  reg  valid_0_11; // @[dcache.scala 93:26]
  reg  valid_0_12; // @[dcache.scala 93:26]
  reg  valid_0_13; // @[dcache.scala 93:26]
  reg  valid_0_14; // @[dcache.scala 93:26]
  reg  valid_0_15; // @[dcache.scala 93:26]
  reg  valid_1_0; // @[dcache.scala 93:26]
  reg  valid_1_1; // @[dcache.scala 93:26]
  reg  valid_1_2; // @[dcache.scala 93:26]
  reg  valid_1_3; // @[dcache.scala 93:26]
  reg  valid_1_4; // @[dcache.scala 93:26]
  reg  valid_1_5; // @[dcache.scala 93:26]
  reg  valid_1_6; // @[dcache.scala 93:26]
  reg  valid_1_7; // @[dcache.scala 93:26]
  reg  valid_1_8; // @[dcache.scala 93:26]
  reg  valid_1_9; // @[dcache.scala 93:26]
  reg  valid_1_10; // @[dcache.scala 93:26]
  reg  valid_1_11; // @[dcache.scala 93:26]
  reg  valid_1_12; // @[dcache.scala 93:26]
  reg  valid_1_13; // @[dcache.scala 93:26]
  reg  valid_1_14; // @[dcache.scala 93:26]
  reg  valid_1_15; // @[dcache.scala 93:26]
  reg  valid_2_0; // @[dcache.scala 93:26]
  reg  valid_2_1; // @[dcache.scala 93:26]
  reg  valid_2_2; // @[dcache.scala 93:26]
  reg  valid_2_3; // @[dcache.scala 93:26]
  reg  valid_2_4; // @[dcache.scala 93:26]
  reg  valid_2_5; // @[dcache.scala 93:26]
  reg  valid_2_6; // @[dcache.scala 93:26]
  reg  valid_2_7; // @[dcache.scala 93:26]
  reg  valid_2_8; // @[dcache.scala 93:26]
  reg  valid_2_9; // @[dcache.scala 93:26]
  reg  valid_2_10; // @[dcache.scala 93:26]
  reg  valid_2_11; // @[dcache.scala 93:26]
  reg  valid_2_12; // @[dcache.scala 93:26]
  reg  valid_2_13; // @[dcache.scala 93:26]
  reg  valid_2_14; // @[dcache.scala 93:26]
  reg  valid_2_15; // @[dcache.scala 93:26]
  reg  valid_3_0; // @[dcache.scala 93:26]
  reg  valid_3_1; // @[dcache.scala 93:26]
  reg  valid_3_2; // @[dcache.scala 93:26]
  reg  valid_3_3; // @[dcache.scala 93:26]
  reg  valid_3_4; // @[dcache.scala 93:26]
  reg  valid_3_5; // @[dcache.scala 93:26]
  reg  valid_3_6; // @[dcache.scala 93:26]
  reg  valid_3_7; // @[dcache.scala 93:26]
  reg  valid_3_8; // @[dcache.scala 93:26]
  reg  valid_3_9; // @[dcache.scala 93:26]
  reg  valid_3_10; // @[dcache.scala 93:26]
  reg  valid_3_11; // @[dcache.scala 93:26]
  reg  valid_3_12; // @[dcache.scala 93:26]
  reg  valid_3_13; // @[dcache.scala 93:26]
  reg  valid_3_14; // @[dcache.scala 93:26]
  reg  valid_3_15; // @[dcache.scala 93:26]
  reg  dirty_0_0; // @[dcache.scala 94:26]
  reg  dirty_0_1; // @[dcache.scala 94:26]
  reg  dirty_0_2; // @[dcache.scala 94:26]
  reg  dirty_0_3; // @[dcache.scala 94:26]
  reg  dirty_0_4; // @[dcache.scala 94:26]
  reg  dirty_0_5; // @[dcache.scala 94:26]
  reg  dirty_0_6; // @[dcache.scala 94:26]
  reg  dirty_0_7; // @[dcache.scala 94:26]
  reg  dirty_0_8; // @[dcache.scala 94:26]
  reg  dirty_0_9; // @[dcache.scala 94:26]
  reg  dirty_0_10; // @[dcache.scala 94:26]
  reg  dirty_0_11; // @[dcache.scala 94:26]
  reg  dirty_0_12; // @[dcache.scala 94:26]
  reg  dirty_0_13; // @[dcache.scala 94:26]
  reg  dirty_0_14; // @[dcache.scala 94:26]
  reg  dirty_0_15; // @[dcache.scala 94:26]
  reg  dirty_1_0; // @[dcache.scala 94:26]
  reg  dirty_1_1; // @[dcache.scala 94:26]
  reg  dirty_1_2; // @[dcache.scala 94:26]
  reg  dirty_1_3; // @[dcache.scala 94:26]
  reg  dirty_1_4; // @[dcache.scala 94:26]
  reg  dirty_1_5; // @[dcache.scala 94:26]
  reg  dirty_1_6; // @[dcache.scala 94:26]
  reg  dirty_1_7; // @[dcache.scala 94:26]
  reg  dirty_1_8; // @[dcache.scala 94:26]
  reg  dirty_1_9; // @[dcache.scala 94:26]
  reg  dirty_1_10; // @[dcache.scala 94:26]
  reg  dirty_1_11; // @[dcache.scala 94:26]
  reg  dirty_1_12; // @[dcache.scala 94:26]
  reg  dirty_1_13; // @[dcache.scala 94:26]
  reg  dirty_1_14; // @[dcache.scala 94:26]
  reg  dirty_1_15; // @[dcache.scala 94:26]
  reg  dirty_2_0; // @[dcache.scala 94:26]
  reg  dirty_2_1; // @[dcache.scala 94:26]
  reg  dirty_2_2; // @[dcache.scala 94:26]
  reg  dirty_2_3; // @[dcache.scala 94:26]
  reg  dirty_2_4; // @[dcache.scala 94:26]
  reg  dirty_2_5; // @[dcache.scala 94:26]
  reg  dirty_2_6; // @[dcache.scala 94:26]
  reg  dirty_2_7; // @[dcache.scala 94:26]
  reg  dirty_2_8; // @[dcache.scala 94:26]
  reg  dirty_2_9; // @[dcache.scala 94:26]
  reg  dirty_2_10; // @[dcache.scala 94:26]
  reg  dirty_2_11; // @[dcache.scala 94:26]
  reg  dirty_2_12; // @[dcache.scala 94:26]
  reg  dirty_2_13; // @[dcache.scala 94:26]
  reg  dirty_2_14; // @[dcache.scala 94:26]
  reg  dirty_2_15; // @[dcache.scala 94:26]
  reg  dirty_3_0; // @[dcache.scala 94:26]
  reg  dirty_3_1; // @[dcache.scala 94:26]
  reg  dirty_3_2; // @[dcache.scala 94:26]
  reg  dirty_3_3; // @[dcache.scala 94:26]
  reg  dirty_3_4; // @[dcache.scala 94:26]
  reg  dirty_3_5; // @[dcache.scala 94:26]
  reg  dirty_3_6; // @[dcache.scala 94:26]
  reg  dirty_3_7; // @[dcache.scala 94:26]
  reg  dirty_3_8; // @[dcache.scala 94:26]
  reg  dirty_3_9; // @[dcache.scala 94:26]
  reg  dirty_3_10; // @[dcache.scala 94:26]
  reg  dirty_3_11; // @[dcache.scala 94:26]
  reg  dirty_3_12; // @[dcache.scala 94:26]
  reg  dirty_3_13; // @[dcache.scala 94:26]
  reg  dirty_3_14; // @[dcache.scala 94:26]
  reg  dirty_3_15; // @[dcache.scala 94:26]
  reg  wait_r; // @[dcache.scala 96:30]
  reg  valid_r; // @[dcache.scala 97:30]
  reg  flush_r; // @[dcache.scala 98:30]
  reg [4:0] mode_r; // @[dcache.scala 99:30]
  reg [63:0] wdata_r; // @[dcache.scala 100:30]
  reg [4:0] amo_r; // @[dcache.scala 101:30]
  wire  _valid_in_T = io_dcRW_dc_mode != 5'h0; // @[dcache.scala 103:40]
  wire  valid_in = io_dcRW_dc_mode != 5'h0 & ~io_flush; // @[dcache.scala 103:54]
  wire  hs_in = _valid_in_T & io_dcRW_ready; // @[dcache.scala 104:52]
  wire  _io_dcRW_ready_T = ~wait_r; // @[dcache.scala 105:34]
  reg [31:0] addr_r; // @[dcache.scala 108:34]
  wire [31:0] cur_addr = hs_in ? io_dcRW_addr : addr_r; // @[dcache.scala 109:30]
  reg [1:0] matchWay_r; // @[dcache.scala 110:34]
  reg [2:0] offset; // @[dcache.scala 111:34]
  reg [63:0] rdatabuf; // @[dcache.scala 112:34]
  wire [3:0] blockIdx = cur_addr[9:6]; // @[dcache.scala 113:35]
  reg [3:0] blockIdx_r; // @[dcache.scala 114:34]
  wire [21:0] cur_tag = cur_addr[31:10]; // @[dcache.scala 115:35]
  wire [21:0] _GEN_1 = 4'h1 == blockIdx ? tag_0_1 : tag_0_0; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_2 = 4'h2 == blockIdx ? tag_0_2 : _GEN_1; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_3 = 4'h3 == blockIdx ? tag_0_3 : _GEN_2; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_4 = 4'h4 == blockIdx ? tag_0_4 : _GEN_3; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_5 = 4'h5 == blockIdx ? tag_0_5 : _GEN_4; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_6 = 4'h6 == blockIdx ? tag_0_6 : _GEN_5; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_7 = 4'h7 == blockIdx ? tag_0_7 : _GEN_6; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_8 = 4'h8 == blockIdx ? tag_0_8 : _GEN_7; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_9 = 4'h9 == blockIdx ? tag_0_9 : _GEN_8; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_10 = 4'ha == blockIdx ? tag_0_10 : _GEN_9; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_11 = 4'hb == blockIdx ? tag_0_11 : _GEN_10; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_12 = 4'hc == blockIdx ? tag_0_12 : _GEN_11; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_13 = 4'hd == blockIdx ? tag_0_13 : _GEN_12; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_14 = 4'he == blockIdx ? tag_0_14 : _GEN_13; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_15 = 4'hf == blockIdx ? tag_0_15 : _GEN_14; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire  _GEN_17 = 4'h1 == blockIdx ? valid_0_1 : valid_0_0; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_18 = 4'h2 == blockIdx ? valid_0_2 : _GEN_17; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_19 = 4'h3 == blockIdx ? valid_0_3 : _GEN_18; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_20 = 4'h4 == blockIdx ? valid_0_4 : _GEN_19; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_21 = 4'h5 == blockIdx ? valid_0_5 : _GEN_20; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_22 = 4'h6 == blockIdx ? valid_0_6 : _GEN_21; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_23 = 4'h7 == blockIdx ? valid_0_7 : _GEN_22; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_24 = 4'h8 == blockIdx ? valid_0_8 : _GEN_23; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_25 = 4'h9 == blockIdx ? valid_0_9 : _GEN_24; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_26 = 4'ha == blockIdx ? valid_0_10 : _GEN_25; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_27 = 4'hb == blockIdx ? valid_0_11 : _GEN_26; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_28 = 4'hc == blockIdx ? valid_0_12 : _GEN_27; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_29 = 4'hd == blockIdx ? valid_0_13 : _GEN_28; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_30 = 4'he == blockIdx ? valid_0_14 : _GEN_29; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_31 = 4'hf == blockIdx ? valid_0_15 : _GEN_30; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  cache_hit_vec_0 = _GEN_15 == cur_tag & _GEN_31; // @[dcache.scala 116:97]
  wire [21:0] _GEN_33 = 4'h1 == blockIdx ? tag_1_1 : tag_1_0; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_34 = 4'h2 == blockIdx ? tag_1_2 : _GEN_33; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_35 = 4'h3 == blockIdx ? tag_1_3 : _GEN_34; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_36 = 4'h4 == blockIdx ? tag_1_4 : _GEN_35; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_37 = 4'h5 == blockIdx ? tag_1_5 : _GEN_36; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_38 = 4'h6 == blockIdx ? tag_1_6 : _GEN_37; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_39 = 4'h7 == blockIdx ? tag_1_7 : _GEN_38; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_40 = 4'h8 == blockIdx ? tag_1_8 : _GEN_39; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_41 = 4'h9 == blockIdx ? tag_1_9 : _GEN_40; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_42 = 4'ha == blockIdx ? tag_1_10 : _GEN_41; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_43 = 4'hb == blockIdx ? tag_1_11 : _GEN_42; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_44 = 4'hc == blockIdx ? tag_1_12 : _GEN_43; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_45 = 4'hd == blockIdx ? tag_1_13 : _GEN_44; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_46 = 4'he == blockIdx ? tag_1_14 : _GEN_45; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_47 = 4'hf == blockIdx ? tag_1_15 : _GEN_46; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire  _GEN_49 = 4'h1 == blockIdx ? valid_1_1 : valid_1_0; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_50 = 4'h2 == blockIdx ? valid_1_2 : _GEN_49; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_51 = 4'h3 == blockIdx ? valid_1_3 : _GEN_50; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_52 = 4'h4 == blockIdx ? valid_1_4 : _GEN_51; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_53 = 4'h5 == blockIdx ? valid_1_5 : _GEN_52; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_54 = 4'h6 == blockIdx ? valid_1_6 : _GEN_53; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_55 = 4'h7 == blockIdx ? valid_1_7 : _GEN_54; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_56 = 4'h8 == blockIdx ? valid_1_8 : _GEN_55; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_57 = 4'h9 == blockIdx ? valid_1_9 : _GEN_56; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_58 = 4'ha == blockIdx ? valid_1_10 : _GEN_57; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_59 = 4'hb == blockIdx ? valid_1_11 : _GEN_58; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_60 = 4'hc == blockIdx ? valid_1_12 : _GEN_59; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_61 = 4'hd == blockIdx ? valid_1_13 : _GEN_60; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_62 = 4'he == blockIdx ? valid_1_14 : _GEN_61; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_63 = 4'hf == blockIdx ? valid_1_15 : _GEN_62; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  cache_hit_vec_1 = _GEN_47 == cur_tag & _GEN_63; // @[dcache.scala 116:97]
  wire [21:0] _GEN_65 = 4'h1 == blockIdx ? tag_2_1 : tag_2_0; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_66 = 4'h2 == blockIdx ? tag_2_2 : _GEN_65; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_67 = 4'h3 == blockIdx ? tag_2_3 : _GEN_66; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_68 = 4'h4 == blockIdx ? tag_2_4 : _GEN_67; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_69 = 4'h5 == blockIdx ? tag_2_5 : _GEN_68; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_70 = 4'h6 == blockIdx ? tag_2_6 : _GEN_69; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_71 = 4'h7 == blockIdx ? tag_2_7 : _GEN_70; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_72 = 4'h8 == blockIdx ? tag_2_8 : _GEN_71; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_73 = 4'h9 == blockIdx ? tag_2_9 : _GEN_72; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_74 = 4'ha == blockIdx ? tag_2_10 : _GEN_73; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_75 = 4'hb == blockIdx ? tag_2_11 : _GEN_74; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_76 = 4'hc == blockIdx ? tag_2_12 : _GEN_75; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_77 = 4'hd == blockIdx ? tag_2_13 : _GEN_76; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_78 = 4'he == blockIdx ? tag_2_14 : _GEN_77; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_79 = 4'hf == blockIdx ? tag_2_15 : _GEN_78; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire  _GEN_81 = 4'h1 == blockIdx ? valid_2_1 : valid_2_0; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_82 = 4'h2 == blockIdx ? valid_2_2 : _GEN_81; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_83 = 4'h3 == blockIdx ? valid_2_3 : _GEN_82; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_84 = 4'h4 == blockIdx ? valid_2_4 : _GEN_83; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_85 = 4'h5 == blockIdx ? valid_2_5 : _GEN_84; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_86 = 4'h6 == blockIdx ? valid_2_6 : _GEN_85; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_87 = 4'h7 == blockIdx ? valid_2_7 : _GEN_86; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_88 = 4'h8 == blockIdx ? valid_2_8 : _GEN_87; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_89 = 4'h9 == blockIdx ? valid_2_9 : _GEN_88; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_90 = 4'ha == blockIdx ? valid_2_10 : _GEN_89; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_91 = 4'hb == blockIdx ? valid_2_11 : _GEN_90; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_92 = 4'hc == blockIdx ? valid_2_12 : _GEN_91; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_93 = 4'hd == blockIdx ? valid_2_13 : _GEN_92; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_94 = 4'he == blockIdx ? valid_2_14 : _GEN_93; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_95 = 4'hf == blockIdx ? valid_2_15 : _GEN_94; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  cache_hit_vec_2 = _GEN_79 == cur_tag & _GEN_95; // @[dcache.scala 116:97]
  wire [21:0] _GEN_97 = 4'h1 == blockIdx ? tag_3_1 : tag_3_0; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_98 = 4'h2 == blockIdx ? tag_3_2 : _GEN_97; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_99 = 4'h3 == blockIdx ? tag_3_3 : _GEN_98; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_100 = 4'h4 == blockIdx ? tag_3_4 : _GEN_99; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_101 = 4'h5 == blockIdx ? tag_3_5 : _GEN_100; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_102 = 4'h6 == blockIdx ? tag_3_6 : _GEN_101; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_103 = 4'h7 == blockIdx ? tag_3_7 : _GEN_102; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_104 = 4'h8 == blockIdx ? tag_3_8 : _GEN_103; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_105 = 4'h9 == blockIdx ? tag_3_9 : _GEN_104; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_106 = 4'ha == blockIdx ? tag_3_10 : _GEN_105; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_107 = 4'hb == blockIdx ? tag_3_11 : _GEN_106; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_108 = 4'hc == blockIdx ? tag_3_12 : _GEN_107; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_109 = 4'hd == blockIdx ? tag_3_13 : _GEN_108; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_110 = 4'he == blockIdx ? tag_3_14 : _GEN_109; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire [21:0] _GEN_111 = 4'hf == blockIdx ? tag_3_15 : _GEN_110; // @[dcache.scala 116:85 dcache.scala 116:85]
  wire  _GEN_113 = 4'h1 == blockIdx ? valid_3_1 : valid_3_0; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_114 = 4'h2 == blockIdx ? valid_3_2 : _GEN_113; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_115 = 4'h3 == blockIdx ? valid_3_3 : _GEN_114; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_116 = 4'h4 == blockIdx ? valid_3_4 : _GEN_115; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_117 = 4'h5 == blockIdx ? valid_3_5 : _GEN_116; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_118 = 4'h6 == blockIdx ? valid_3_6 : _GEN_117; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_119 = 4'h7 == blockIdx ? valid_3_7 : _GEN_118; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_120 = 4'h8 == blockIdx ? valid_3_8 : _GEN_119; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_121 = 4'h9 == blockIdx ? valid_3_9 : _GEN_120; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_122 = 4'ha == blockIdx ? valid_3_10 : _GEN_121; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_123 = 4'hb == blockIdx ? valid_3_11 : _GEN_122; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_124 = 4'hc == blockIdx ? valid_3_12 : _GEN_123; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_125 = 4'hd == blockIdx ? valid_3_13 : _GEN_124; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_126 = 4'he == blockIdx ? valid_3_14 : _GEN_125; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  _GEN_127 = 4'hf == blockIdx ? valid_3_15 : _GEN_126; // @[dcache.scala 116:97 dcache.scala 116:97]
  wire  cache_hit_vec_3 = _GEN_111 == cur_tag & _GEN_127; // @[dcache.scala 116:97]
  wire [3:0] _cacheHit_T = {cache_hit_vec_3,cache_hit_vec_2,cache_hit_vec_1,cache_hit_vec_0}; // @[dcache.scala 117:47]
  wire  cacheHit = |_cacheHit_T; // @[dcache.scala 117:50]
  wire [1:0] matchWay_hi_1 = _cacheHit_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] matchWay_lo_1 = _cacheHit_T[1:0]; // @[OneHot.scala 31:18]
  wire  matchWay_hi_2 = |matchWay_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _matchWay_T_1 = matchWay_hi_1 | matchWay_lo_1; // @[OneHot.scala 32:28]
  wire  matchWay_lo_2 = _matchWay_T_1[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] _matchWay_T_2 = {matchWay_hi_2,matchWay_lo_2}; // @[Cat.scala 30:58]
  wire [2:0] _matchWay_T_3 = {matchWay_prng_io_out_2,matchWay_prng_io_out_1,matchWay_prng_io_out_0}; // @[PRNG.scala 86:17]
  wire [1:0] _matchWay_T_5 = hs_in ? _matchWay_T_3[2:1] : matchWay_r; // @[dcache.scala 118:69]
  wire [1:0] matchWay = cacheHit ? _matchWay_T_2 : _matchWay_T_5; // @[dcache.scala 118:30]
  wire [1:0] _GEN_129 = hs_in ? matchWay : matchWay_r; // @[dcache.scala 120:16 dcache.scala 122:20 dcache.scala 110:34]
  wire [4:0] _GEN_130 = hs_in ? io_dcRW_dc_mode : mode_r; // @[dcache.scala 120:16 dcache.scala 123:17 dcache.scala 99:30]
  wire [63:0] _GEN_131 = hs_in ? io_dcRW_wdata : wdata_r; // @[dcache.scala 120:16 dcache.scala 124:17 dcache.scala 100:30]
  wire [3:0] _GEN_133 = hs_in ? io_dcRW_addr[9:6] : blockIdx_r; // @[dcache.scala 120:16 dcache.scala 126:20 dcache.scala 114:34]
  wire  _GEN_134 = io_flush | flush_r; // @[dcache.scala 129:19 dcache.scala 130:17 dcache.scala 98:30]
  wire  _GEN_136 = valid_0_0 & dirty_0_0 ? 1'h0 : 1'h1; // @[dcache.scala 138:45 dcache.scala 141:28 dcache.scala 135:52]
  wire  _T_1 = valid_0_1 & dirty_0_1; // @[dcache.scala 138:30]
  wire  _GEN_139 = valid_0_1 & dirty_0_1 ? 1'h0 : _GEN_136; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_141 = valid_0_2 & dirty_0_2 ? 2'h2 : {{1'd0}, _T_1}; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_142 = valid_0_2 & dirty_0_2 ? 1'h0 : _GEN_139; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_144 = valid_0_3 & dirty_0_3 ? 2'h3 : _GEN_141; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_145 = valid_0_3 & dirty_0_3 ? 1'h0 : _GEN_142; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [2:0] _GEN_147 = valid_0_4 & dirty_0_4 ? 3'h4 : {{1'd0}, _GEN_144}; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_148 = valid_0_4 & dirty_0_4 ? 1'h0 : _GEN_145; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [2:0] _GEN_150 = valid_0_5 & dirty_0_5 ? 3'h5 : _GEN_147; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_151 = valid_0_5 & dirty_0_5 ? 1'h0 : _GEN_148; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [2:0] _GEN_153 = valid_0_6 & dirty_0_6 ? 3'h6 : _GEN_150; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_154 = valid_0_6 & dirty_0_6 ? 1'h0 : _GEN_151; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [2:0] _GEN_156 = valid_0_7 & dirty_0_7 ? 3'h7 : _GEN_153; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_157 = valid_0_7 & dirty_0_7 ? 1'h0 : _GEN_154; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_159 = valid_0_8 & dirty_0_8 ? 4'h8 : {{1'd0}, _GEN_156}; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_160 = valid_0_8 & dirty_0_8 ? 1'h0 : _GEN_157; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_162 = valid_0_9 & dirty_0_9 ? 4'h9 : _GEN_159; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_163 = valid_0_9 & dirty_0_9 ? 1'h0 : _GEN_160; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_165 = valid_0_10 & dirty_0_10 ? 4'ha : _GEN_162; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_166 = valid_0_10 & dirty_0_10 ? 1'h0 : _GEN_163; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_168 = valid_0_11 & dirty_0_11 ? 4'hb : _GEN_165; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_169 = valid_0_11 & dirty_0_11 ? 1'h0 : _GEN_166; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_171 = valid_0_12 & dirty_0_12 ? 4'hc : _GEN_168; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_172 = valid_0_12 & dirty_0_12 ? 1'h0 : _GEN_169; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_174 = valid_0_13 & dirty_0_13 ? 4'hd : _GEN_171; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_175 = valid_0_13 & dirty_0_13 ? 1'h0 : _GEN_172; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_177 = valid_0_14 & dirty_0_14 ? 4'he : _GEN_174; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_178 = valid_0_14 & dirty_0_14 ? 1'h0 : _GEN_175; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_180 = valid_0_15 & dirty_0_15 ? 4'hf : _GEN_177; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_181 = valid_0_15 & dirty_0_15 ? 1'h0 : _GEN_178; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_183 = valid_1_0 & dirty_1_0 ? 4'h0 : _GEN_180; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_184 = valid_1_0 & dirty_1_0 ? 1'h0 : _GEN_181; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_186 = valid_1_1 & dirty_1_1 ? 4'h1 : _GEN_183; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_187 = valid_1_1 & dirty_1_1 ? 1'h0 : _GEN_184; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_189 = valid_1_2 & dirty_1_2 ? 4'h2 : _GEN_186; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_190 = valid_1_2 & dirty_1_2 ? 1'h0 : _GEN_187; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_192 = valid_1_3 & dirty_1_3 ? 4'h3 : _GEN_189; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_193 = valid_1_3 & dirty_1_3 ? 1'h0 : _GEN_190; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_195 = valid_1_4 & dirty_1_4 ? 4'h4 : _GEN_192; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_196 = valid_1_4 & dirty_1_4 ? 1'h0 : _GEN_193; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_198 = valid_1_5 & dirty_1_5 ? 4'h5 : _GEN_195; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_199 = valid_1_5 & dirty_1_5 ? 1'h0 : _GEN_196; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_201 = valid_1_6 & dirty_1_6 ? 4'h6 : _GEN_198; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_202 = valid_1_6 & dirty_1_6 ? 1'h0 : _GEN_199; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_204 = valid_1_7 & dirty_1_7 ? 4'h7 : _GEN_201; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_205 = valid_1_7 & dirty_1_7 ? 1'h0 : _GEN_202; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_207 = valid_1_8 & dirty_1_8 ? 4'h8 : _GEN_204; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_208 = valid_1_8 & dirty_1_8 ? 1'h0 : _GEN_205; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_210 = valid_1_9 & dirty_1_9 ? 4'h9 : _GEN_207; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_211 = valid_1_9 & dirty_1_9 ? 1'h0 : _GEN_208; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_213 = valid_1_10 & dirty_1_10 ? 4'ha : _GEN_210; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_214 = valid_1_10 & dirty_1_10 ? 1'h0 : _GEN_211; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_216 = valid_1_11 & dirty_1_11 ? 4'hb : _GEN_213; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_217 = valid_1_11 & dirty_1_11 ? 1'h0 : _GEN_214; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_219 = valid_1_12 & dirty_1_12 ? 4'hc : _GEN_216; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_220 = valid_1_12 & dirty_1_12 ? 1'h0 : _GEN_217; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [3:0] _GEN_222 = valid_1_13 & dirty_1_13 ? 4'hd : _GEN_219; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_223 = valid_1_13 & dirty_1_13 ? 1'h0 : _GEN_220; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire  _GEN_224 = valid_1_14 & dirty_1_14 | (valid_1_13 & dirty_1_13 | (valid_1_12 & dirty_1_12 | (valid_1_11 &
    dirty_1_11 | (valid_1_10 & dirty_1_10 | (valid_1_9 & dirty_1_9 | (valid_1_8 & dirty_1_8 | (valid_1_7 & dirty_1_7 | (
    valid_1_6 & dirty_1_6 | (valid_1_5 & dirty_1_5 | (valid_1_4 & dirty_1_4 | (valid_1_3 & dirty_1_3 | (valid_1_2 &
    dirty_1_2 | (valid_1_1 & dirty_1_1 | valid_1_0 & dirty_1_0))))))))))))); // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_225 = valid_1_14 & dirty_1_14 ? 4'he : _GEN_222; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_226 = valid_1_14 & dirty_1_14 ? 1'h0 : _GEN_223; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire  _GEN_227 = valid_1_15 & dirty_1_15 | _GEN_224; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_228 = valid_1_15 & dirty_1_15 ? 4'hf : _GEN_225; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_229 = valid_1_15 & dirty_1_15 ? 1'h0 : _GEN_226; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_230 = valid_2_0 & dirty_2_0 ? 2'h2 : {{1'd0}, _GEN_227}; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_231 = valid_2_0 & dirty_2_0 ? 4'h0 : _GEN_228; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_232 = valid_2_0 & dirty_2_0 ? 1'h0 : _GEN_229; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_233 = valid_2_1 & dirty_2_1 ? 2'h2 : _GEN_230; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_234 = valid_2_1 & dirty_2_1 ? 4'h1 : _GEN_231; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_235 = valid_2_1 & dirty_2_1 ? 1'h0 : _GEN_232; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_236 = valid_2_2 & dirty_2_2 ? 2'h2 : _GEN_233; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_237 = valid_2_2 & dirty_2_2 ? 4'h2 : _GEN_234; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_238 = valid_2_2 & dirty_2_2 ? 1'h0 : _GEN_235; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_239 = valid_2_3 & dirty_2_3 ? 2'h2 : _GEN_236; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_240 = valid_2_3 & dirty_2_3 ? 4'h3 : _GEN_237; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_241 = valid_2_3 & dirty_2_3 ? 1'h0 : _GEN_238; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_242 = valid_2_4 & dirty_2_4 ? 2'h2 : _GEN_239; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_243 = valid_2_4 & dirty_2_4 ? 4'h4 : _GEN_240; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_244 = valid_2_4 & dirty_2_4 ? 1'h0 : _GEN_241; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_245 = valid_2_5 & dirty_2_5 ? 2'h2 : _GEN_242; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_246 = valid_2_5 & dirty_2_5 ? 4'h5 : _GEN_243; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_247 = valid_2_5 & dirty_2_5 ? 1'h0 : _GEN_244; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_248 = valid_2_6 & dirty_2_6 ? 2'h2 : _GEN_245; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_249 = valid_2_6 & dirty_2_6 ? 4'h6 : _GEN_246; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_250 = valid_2_6 & dirty_2_6 ? 1'h0 : _GEN_247; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_251 = valid_2_7 & dirty_2_7 ? 2'h2 : _GEN_248; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_252 = valid_2_7 & dirty_2_7 ? 4'h7 : _GEN_249; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_253 = valid_2_7 & dirty_2_7 ? 1'h0 : _GEN_250; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_254 = valid_2_8 & dirty_2_8 ? 2'h2 : _GEN_251; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_255 = valid_2_8 & dirty_2_8 ? 4'h8 : _GEN_252; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_256 = valid_2_8 & dirty_2_8 ? 1'h0 : _GEN_253; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_257 = valid_2_9 & dirty_2_9 ? 2'h2 : _GEN_254; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_258 = valid_2_9 & dirty_2_9 ? 4'h9 : _GEN_255; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_259 = valid_2_9 & dirty_2_9 ? 1'h0 : _GEN_256; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_260 = valid_2_10 & dirty_2_10 ? 2'h2 : _GEN_257; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_261 = valid_2_10 & dirty_2_10 ? 4'ha : _GEN_258; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_262 = valid_2_10 & dirty_2_10 ? 1'h0 : _GEN_259; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_263 = valid_2_11 & dirty_2_11 ? 2'h2 : _GEN_260; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_264 = valid_2_11 & dirty_2_11 ? 4'hb : _GEN_261; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_265 = valid_2_11 & dirty_2_11 ? 1'h0 : _GEN_262; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_266 = valid_2_12 & dirty_2_12 ? 2'h2 : _GEN_263; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_267 = valid_2_12 & dirty_2_12 ? 4'hc : _GEN_264; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_268 = valid_2_12 & dirty_2_12 ? 1'h0 : _GEN_265; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_269 = valid_2_13 & dirty_2_13 ? 2'h2 : _GEN_266; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_270 = valid_2_13 & dirty_2_13 ? 4'hd : _GEN_267; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_271 = valid_2_13 & dirty_2_13 ? 1'h0 : _GEN_268; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_272 = valid_2_14 & dirty_2_14 ? 2'h2 : _GEN_269; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_273 = valid_2_14 & dirty_2_14 ? 4'he : _GEN_270; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_274 = valid_2_14 & dirty_2_14 ? 1'h0 : _GEN_271; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_275 = valid_2_15 & dirty_2_15 ? 2'h2 : _GEN_272; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_276 = valid_2_15 & dirty_2_15 ? 4'hf : _GEN_273; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_277 = valid_2_15 & dirty_2_15 ? 1'h0 : _GEN_274; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_278 = valid_3_0 & dirty_3_0 ? 2'h3 : _GEN_275; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_279 = valid_3_0 & dirty_3_0 ? 4'h0 : _GEN_276; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_280 = valid_3_0 & dirty_3_0 ? 1'h0 : _GEN_277; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_281 = valid_3_1 & dirty_3_1 ? 2'h3 : _GEN_278; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_282 = valid_3_1 & dirty_3_1 ? 4'h1 : _GEN_279; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_283 = valid_3_1 & dirty_3_1 ? 1'h0 : _GEN_280; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_284 = valid_3_2 & dirty_3_2 ? 2'h3 : _GEN_281; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_285 = valid_3_2 & dirty_3_2 ? 4'h2 : _GEN_282; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_286 = valid_3_2 & dirty_3_2 ? 1'h0 : _GEN_283; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_287 = valid_3_3 & dirty_3_3 ? 2'h3 : _GEN_284; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_288 = valid_3_3 & dirty_3_3 ? 4'h3 : _GEN_285; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_289 = valid_3_3 & dirty_3_3 ? 1'h0 : _GEN_286; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_290 = valid_3_4 & dirty_3_4 ? 2'h3 : _GEN_287; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_291 = valid_3_4 & dirty_3_4 ? 4'h4 : _GEN_288; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_292 = valid_3_4 & dirty_3_4 ? 1'h0 : _GEN_289; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_293 = valid_3_5 & dirty_3_5 ? 2'h3 : _GEN_290; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_294 = valid_3_5 & dirty_3_5 ? 4'h5 : _GEN_291; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_295 = valid_3_5 & dirty_3_5 ? 1'h0 : _GEN_292; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_296 = valid_3_6 & dirty_3_6 ? 2'h3 : _GEN_293; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_297 = valid_3_6 & dirty_3_6 ? 4'h6 : _GEN_294; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_298 = valid_3_6 & dirty_3_6 ? 1'h0 : _GEN_295; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_299 = valid_3_7 & dirty_3_7 ? 2'h3 : _GEN_296; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_300 = valid_3_7 & dirty_3_7 ? 4'h7 : _GEN_297; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_301 = valid_3_7 & dirty_3_7 ? 1'h0 : _GEN_298; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_302 = valid_3_8 & dirty_3_8 ? 2'h3 : _GEN_299; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_303 = valid_3_8 & dirty_3_8 ? 4'h8 : _GEN_300; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_304 = valid_3_8 & dirty_3_8 ? 1'h0 : _GEN_301; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_305 = valid_3_9 & dirty_3_9 ? 2'h3 : _GEN_302; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_306 = valid_3_9 & dirty_3_9 ? 4'h9 : _GEN_303; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_307 = valid_3_9 & dirty_3_9 ? 1'h0 : _GEN_304; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_308 = valid_3_10 & dirty_3_10 ? 2'h3 : _GEN_305; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_309 = valid_3_10 & dirty_3_10 ? 4'ha : _GEN_306; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_310 = valid_3_10 & dirty_3_10 ? 1'h0 : _GEN_307; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_311 = valid_3_11 & dirty_3_11 ? 2'h3 : _GEN_308; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_312 = valid_3_11 & dirty_3_11 ? 4'hb : _GEN_309; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_313 = valid_3_11 & dirty_3_11 ? 1'h0 : _GEN_310; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_314 = valid_3_12 & dirty_3_12 ? 2'h3 : _GEN_311; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_315 = valid_3_12 & dirty_3_12 ? 4'hc : _GEN_312; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_316 = valid_3_12 & dirty_3_12 ? 1'h0 : _GEN_313; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_317 = valid_3_13 & dirty_3_13 ? 2'h3 : _GEN_314; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_318 = valid_3_13 & dirty_3_13 ? 4'hd : _GEN_315; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_319 = valid_3_13 & dirty_3_13 ? 1'h0 : _GEN_316; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] _GEN_320 = valid_3_14 & dirty_3_14 ? 2'h3 : _GEN_317; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] _GEN_321 = valid_3_14 & dirty_3_14 ? 4'he : _GEN_318; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  _GEN_322 = valid_3_14 & dirty_3_14 ? 1'h0 : _GEN_319; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [1:0] flush_way = valid_3_15 & dirty_3_15 ? 2'h3 : _GEN_320; // @[dcache.scala 138:45 dcache.scala 139:27]
  wire [3:0] flush_idx = valid_3_15 & dirty_3_15 ? 4'hf : _GEN_321; // @[dcache.scala 138:45 dcache.scala 140:27]
  wire  flush_done = valid_3_15 & dirty_3_15 ? 1'h0 : _GEN_322; // @[dcache.scala 138:45 dcache.scala 141:28]
  wire [5:0] cur_ram_addr = cur_addr[9:4]; // @[dcache.scala 146:35]
  wire [1:0] cur_axi_addr_lo = offset[2:1]; // @[dcache.scala 147:61]
  wire [5:0] _cur_axi_addr_T = {flush_idx,cur_axi_addr_lo}; // @[Cat.scala 30:58]
  wire [5:0] _cur_axi_addr_T_1 = {blockIdx,cur_axi_addr_lo}; // @[Cat.scala 30:58]
  wire [5:0] cur_axi_addr = flush_r ? _cur_axi_addr_T : _cur_axi_addr_T_1; // @[dcache.scala 147:30]
  wire [3:0] pre_blockIdx = addr_r[9:6]; // @[dcache.scala 150:33]
  wire [21:0] pre_tag = addr_r[31:10]; // @[dcache.scala 151:29]
  reg [2:0] state; // @[dcache.scala 153:24]
  wire  _rdata128_T = 2'h1 == matchWay_r; // @[Mux.scala 80:60]
  wire [127:0] _rdata128_T_1 = 2'h1 == matchWay_r ? io_dc2sr1_rdata : io_dc2sr0_rdata; // @[Mux.scala 80:57]
  wire  _rdata128_T_2 = 2'h2 == matchWay_r; // @[Mux.scala 80:60]
  wire [127:0] _rdata128_T_3 = 2'h2 == matchWay_r ? io_dc2sr2_rdata : _rdata128_T_1; // @[Mux.scala 80:57]
  wire  _rdata128_T_4 = 2'h3 == matchWay_r; // @[Mux.scala 80:60]
  wire [127:0] rdata128 = 2'h3 == matchWay_r ? io_dc2sr3_rdata : _rdata128_T_3; // @[Mux.scala 80:57]
  wire [3:0] rdata64_hi = addr_r[3:0]; // @[dcache.scala 160:41]
  wire [6:0] _rdata64_T = {rdata64_hi,3'h0}; // @[Cat.scala 30:58]
  wire [127:0] rdata64 = rdata128 >> _rdata64_T; // @[dcache.scala 160:28]
  wire [55:0] io_dcRW_rdata_hi = rdata64[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_dcRW_rdata_lo = rdata64[7:0]; // @[common.scala 296:70]
  wire [63:0] _io_dcRW_rdata_T_2 = {io_dcRW_rdata_hi,io_dcRW_rdata_lo}; // @[Cat.scala 30:58]
  wire [47:0] io_dcRW_rdata_hi_1 = rdata64[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [15:0] io_dcRW_rdata_lo_1 = rdata64[15:0]; // @[common.scala 298:72]
  wire [63:0] _io_dcRW_rdata_T_6 = {io_dcRW_rdata_hi_1,io_dcRW_rdata_lo_1}; // @[Cat.scala 30:58]
  wire [31:0] io_dcRW_rdata_hi_2 = rdata64[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] io_dcRW_rdata_lo_2 = rdata64[31:0]; // @[common.scala 300:72]
  wire [63:0] _io_dcRW_rdata_T_10 = {io_dcRW_rdata_hi_2,io_dcRW_rdata_lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _io_dcRW_rdata_T_16 = 5'h4 == mode_r ? _io_dcRW_rdata_T_2 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_dcRW_rdata_T_18 = 5'h14 == mode_r ? {{56'd0}, io_dcRW_rdata_lo} : _io_dcRW_rdata_T_16; // @[Mux.scala 80:57]
  wire [63:0] _io_dcRW_rdata_T_20 = 5'h5 == mode_r ? _io_dcRW_rdata_T_6 : _io_dcRW_rdata_T_18; // @[Mux.scala 80:57]
  wire [63:0] _io_dcRW_rdata_T_22 = 5'h15 == mode_r ? {{48'd0}, io_dcRW_rdata_lo_1} : _io_dcRW_rdata_T_20; // @[Mux.scala 80:57]
  wire [63:0] _io_dcRW_rdata_T_24 = 5'h6 == mode_r ? _io_dcRW_rdata_T_10 : _io_dcRW_rdata_T_22; // @[Mux.scala 80:57]
  wire [63:0] _io_dcRW_rdata_T_26 = 5'h16 == mode_r ? {{32'd0}, io_dcRW_rdata_lo_2} : _io_dcRW_rdata_T_24; // @[Mux.scala 80:57]
  wire [127:0] _io_dcRW_rdata_T_28 = 5'h7 == mode_r ? rdata64 : {{64'd0}, _io_dcRW_rdata_T_26}; // @[Mux.scala 80:57]
  wire [127:0] _io_dcRW_rdata_T_30 = 5'he == mode_r ? {{64'd0}, _io_dcRW_rdata_T_10} : _io_dcRW_rdata_T_28; // @[Mux.scala 80:57]
  wire [127:0] _io_dcRW_rdata_T_32 = 5'hf == mode_r ? rdata64 : _io_dcRW_rdata_T_30; // @[Mux.scala 80:57]
  wire [1:0] cur_mode_sl = _GEN_130[3:2]; // @[dcache.scala 162:31]
  wire  cur_mode_s = _GEN_130[3]; // @[dcache.scala 163:31]
  wire [63:0] _amo_rdata_ans_T_11 = 2'h2 == mode_r[1:0] ? _io_dcRW_rdata_T_10 : rdata64[63:0]; // @[Mux.scala 80:57]
  wire [63:0] _amo_rdata_ans_T_13 = 2'h1 == mode_r[1:0] ? _io_dcRW_rdata_T_6 : _amo_rdata_ans_T_11; // @[Mux.scala 80:57]
  wire [63:0] amo_rdata = 2'h0 == mode_r[1:0] ? _io_dcRW_rdata_T_2 : _amo_rdata_ans_T_13; // @[Mux.scala 80:57]
  wire [31:0] amo_imm_ans_hi = wdata_r[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] amo_imm_ans_lo = wdata_r[31:0]; // @[common.scala 319:48]
  wire [63:0] _amo_imm_ans_T_3 = {amo_imm_ans_hi,amo_imm_ans_lo}; // @[Cat.scala 30:58]
  wire [47:0] amo_imm_ans_hi_1 = wdata_r[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [15:0] amo_imm_ans_lo_1 = wdata_r[15:0]; // @[common.scala 320:48]
  wire [63:0] _amo_imm_ans_T_6 = {amo_imm_ans_hi_1,amo_imm_ans_lo_1}; // @[Cat.scala 30:58]
  wire [55:0] amo_imm_ans_hi_2 = wdata_r[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [7:0] amo_imm_ans_lo_2 = wdata_r[7:0]; // @[common.scala 321:47]
  wire [63:0] _amo_imm_ans_T_9 = {amo_imm_ans_hi_2,amo_imm_ans_lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _amo_imm_ans_T_11 = 2'h2 == mode_r[1:0] ? _amo_imm_ans_T_3 : wdata_r; // @[Mux.scala 80:57]
  wire [63:0] _amo_imm_ans_T_13 = 2'h1 == mode_r[1:0] ? _amo_imm_ans_T_6 : _amo_imm_ans_T_11; // @[Mux.scala 80:57]
  wire [63:0] amo_imm = 2'h0 == mode_r[1:0] ? _amo_imm_ans_T_9 : _amo_imm_ans_T_13; // @[Mux.scala 80:57]
  wire [63:0] _amo_alu_T_1 = amo_imm + amo_rdata; // @[dcache.scala 172:29]
  wire [63:0] _amo_alu_T_2 = amo_imm ^ amo_rdata; // @[dcache.scala 173:29]
  wire [63:0] _amo_alu_T_3 = amo_imm & amo_rdata; // @[dcache.scala 174:29]
  wire [63:0] _amo_alu_T_4 = amo_imm | amo_rdata; // @[dcache.scala 175:29]
  wire [63:0] _amo_alu_T_5 = 2'h0 == mode_r[1:0] ? _amo_imm_ans_T_9 : _amo_imm_ans_T_13; // @[dcache.scala 176:32]
  wire [63:0] _amo_alu_T_6 = 2'h0 == mode_r[1:0] ? _io_dcRW_rdata_T_2 : _amo_rdata_ans_T_13; // @[dcache.scala 176:51]
  wire  _amo_alu_T_7 = $signed(_amo_alu_T_5) > $signed(_amo_alu_T_6); // @[dcache.scala 176:39]
  wire [63:0] _amo_alu_T_8 = $signed(_amo_alu_T_5) > $signed(_amo_alu_T_6) ? amo_rdata : amo_imm; // @[dcache.scala 176:23]
  wire [63:0] _amo_alu_T_12 = _amo_alu_T_7 ? amo_imm : amo_rdata; // @[dcache.scala 177:23]
  wire  _amo_alu_T_13 = amo_imm > amo_rdata; // @[dcache.scala 178:32]
  wire [63:0] _amo_alu_T_14 = amo_imm > amo_rdata ? amo_rdata : amo_imm; // @[dcache.scala 178:23]
  wire [63:0] _amo_alu_T_16 = _amo_alu_T_13 ? amo_imm : amo_rdata; // @[dcache.scala 179:23]
  wire [63:0] _amo_alu_T_18 = 5'h1 == amo_r ? amo_imm : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _amo_alu_T_20 = 5'h0 == amo_r ? _amo_alu_T_1 : _amo_alu_T_18; // @[Mux.scala 80:57]
  wire [63:0] _amo_alu_T_22 = 5'h4 == amo_r ? _amo_alu_T_2 : _amo_alu_T_20; // @[Mux.scala 80:57]
  wire [63:0] _amo_alu_T_24 = 5'hc == amo_r ? _amo_alu_T_3 : _amo_alu_T_22; // @[Mux.scala 80:57]
  wire [63:0] _amo_alu_T_26 = 5'h8 == amo_r ? _amo_alu_T_4 : _amo_alu_T_24; // @[Mux.scala 80:57]
  wire [63:0] _amo_alu_T_28 = 5'h10 == amo_r ? _amo_alu_T_8 : _amo_alu_T_26; // @[Mux.scala 80:57]
  wire [63:0] _amo_alu_T_30 = 5'h14 == amo_r ? _amo_alu_T_12 : _amo_alu_T_28; // @[Mux.scala 80:57]
  wire [63:0] _amo_alu_T_32 = 5'h1c == amo_r ? _amo_alu_T_14 : _amo_alu_T_30; // @[Mux.scala 80:57]
  wire [63:0] amo_alu = 5'h1c == amo_r ? _amo_alu_T_16 : _amo_alu_T_32; // @[Mux.scala 80:57]
  wire [31:0] amo_wdata_ans_lo = amo_alu[31:0]; // @[common.scala 310:39]
  wire [63:0] _amo_wdata_ans_T_1 = {32'h0,amo_wdata_ans_lo}; // @[Cat.scala 30:58]
  wire [15:0] amo_wdata_ans_lo_1 = amo_alu[15:0]; // @[common.scala 311:39]
  wire [63:0] _amo_wdata_ans_T_2 = {48'h0,amo_wdata_ans_lo_1}; // @[Cat.scala 30:58]
  wire [7:0] amo_wdata_ans_lo_2 = amo_alu[7:0]; // @[common.scala 312:39]
  wire [63:0] _amo_wdata_ans_T_3 = {56'h0,amo_wdata_ans_lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _amo_wdata_ans_T_5 = 2'h2 == mode_r[1:0] ? _amo_wdata_ans_T_1 : amo_alu; // @[Mux.scala 80:57]
  wire [63:0] _amo_wdata_ans_T_7 = 2'h1 == mode_r[1:0] ? _amo_wdata_ans_T_2 : _amo_wdata_ans_T_5; // @[Mux.scala 80:57]
  wire [63:0] amo_wdata_ans = 2'h0 == mode_r[1:0] ? _amo_wdata_ans_T_3 : _amo_wdata_ans_T_7; // @[Mux.scala 80:57]
  wire [3:0] amo_wdata_hi = cur_addr[3:0]; // @[dcache.scala 181:76]
  wire [6:0] _amo_wdata_T_1 = {amo_wdata_hi,3'h0}; // @[Cat.scala 30:58]
  wire [190:0] _GEN_2500 = {{127'd0}, amo_wdata_ans}; // @[dcache.scala 181:60]
  wire [190:0] amo_wdata = _GEN_2500 << _amo_wdata_T_1; // @[dcache.scala 181:60]
  wire [190:0] _GEN_2501 = {{127'd0}, _GEN_131}; // @[dcache.scala 183:32]
  wire [190:0] inp_wdata = _GEN_2501 << _amo_wdata_T_1; // @[dcache.scala 183:32]
  wire [127:0] _inp_mask_T_2 = 2'h1 == _GEN_130[1:0] ? 128'hffff : 128'hff; // @[Mux.scala 80:57]
  wire [127:0] _inp_mask_T_4 = 2'h2 == _GEN_130[1:0] ? 128'hffffffff : _inp_mask_T_2; // @[Mux.scala 80:57]
  wire [127:0] _inp_mask_T_6 = 2'h3 == _GEN_130[1:0] ? 128'hffffffffffffffff : _inp_mask_T_4; // @[Mux.scala 80:57]
  wire [254:0] _GEN_2502 = {{127'd0}, _inp_mask_T_6}; // @[dcache.scala 189:24]
  wire [254:0] inp_mask = _GEN_2502 << _amo_wdata_T_1; // @[dcache.scala 189:24]
  wire  _io_dc2sr0_addr_T = state == 3'h0; // @[dcache.scala 190:33]
  wire  _io_dc2sr0_addr_T_1 = state == 3'h5; // @[dcache.scala 190:52]
  wire  _io_dc2sr0_addr_T_2 = state == 3'h0 | state == 3'h5; // @[dcache.scala 190:43]
  wire  _io_dc2sr0_cen_T_2 = wait_r | hs_in | flush_r; // @[dcache.scala 194:60]
  wire  _T_68 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_73 = cur_mode_sl == 2'h3; // @[dcache.scala 234:34]
  wire  _GEN_521 = cur_mode_sl == 2'h3 ? 1'h0 : cur_mode_s; // @[dcache.scala 234:42 dcache.scala 211:13 dcache.scala 239:25]
  wire  _GEN_593 = cacheHit & _GEN_521; // @[dcache.scala 233:33 dcache.scala 211:13]
  wire  _GEN_600 = ~hs_in & _io_dcRW_ready_T ? 1'h0 : _GEN_593; // @[dcache.scala 231:42 dcache.scala 211:13]
  wire  _GEN_607 = flush_r | io_flush ? 1'h0 : _GEN_600; // @[dcache.scala 229:38 dcache.scala 211:13]
  wire  _T_74 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_76 = 3'h2 == state; // @[Conditional.scala 37:30]
  reg  axiRdataEn; // @[dcache.scala 220:34]
  wire  _GEN_875 = axiRdataEn & io_dataAxi_rd_valid & offset[0]; // @[dcache.scala 265:52 dcache.scala 211:13]
  wire  _T_79 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_81 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_83 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_1740 = _T_81 ? 1'h0 : _T_83; // @[Conditional.scala 39:67 dcache.scala 211:13]
  wire  _GEN_1879 = _T_79 ? 1'h0 : _GEN_1740; // @[Conditional.scala 39:67 dcache.scala 211:13]
  wire  _GEN_1886 = _T_76 ? _GEN_875 : _GEN_1879; // @[Conditional.scala 39:67]
  wire  _GEN_2093 = _T_74 ? 1'h0 : _GEN_1886; // @[Conditional.scala 39:67 dcache.scala 211:13]
  wire  wen = _T_68 ? _GEN_607 : _GEN_2093; // @[Conditional.scala 40:58]
  wire [127:0] _io_dc2sr0_wdata_T_2 = {io_dataAxi_rd_bits_data,rdatabuf}; // @[Cat.scala 30:58]
  wire [190:0] _io_dc2sr0_wdata_T_3 = _io_dc2sr0_addr_T ? inp_wdata : {{63'd0}, _io_dc2sr0_wdata_T_2}; // @[dcache.scala 203:28]
  wire [190:0] _io_dc2sr0_wdata_T_4 = _io_dc2sr0_addr_T_1 ? amo_wdata : _io_dc2sr0_wdata_T_3; // @[dcache.scala 202:27]
  wire [254:0] _GEN_522 = cur_mode_sl == 2'h3 ? 255'hffffffffffffffffffffffffffffffff : inp_mask; // @[dcache.scala 234:42 dcache.scala 212:13 dcache.scala 240:26]
  wire [254:0] _GEN_594 = cacheHit ? _GEN_522 : 255'hffffffffffffffffffffffffffffffff; // @[dcache.scala 233:33 dcache.scala 212:13]
  wire [254:0] _GEN_601 = ~hs_in & _io_dcRW_ready_T ? 255'hffffffffffffffffffffffffffffffff : _GEN_594; // @[dcache.scala 231:42 dcache.scala 212:13]
  wire [254:0] _GEN_608 = flush_r | io_flush ? 255'hffffffffffffffffffffffffffffffff : _GEN_601; // @[dcache.scala 229:38 dcache.scala 212:13]
  wire [254:0] _GEN_1538 = _T_83 ? inp_mask : 255'hffffffffffffffffffffffffffffffff; // @[Conditional.scala 39:67 dcache.scala 303:21 dcache.scala 212:13]
  wire [254:0] _GEN_1741 = _T_81 ? 255'hffffffffffffffffffffffffffffffff : _GEN_1538; // @[Conditional.scala 39:67 dcache.scala 212:13]
  wire [254:0] _GEN_1880 = _T_79 ? 255'hffffffffffffffffffffffffffffffff : _GEN_1741; // @[Conditional.scala 39:67 dcache.scala 212:13]
  wire [254:0] _GEN_2084 = _T_76 ? 255'hffffffffffffffffffffffffffffffff : _GEN_1880; // @[Conditional.scala 39:67 dcache.scala 212:13]
  wire [254:0] _GEN_2289 = _T_74 ? 255'hffffffffffffffffffffffffffffffff : _GEN_2084; // @[Conditional.scala 39:67 dcache.scala 212:13]
  wire [254:0] _GEN_2298 = _T_68 ? _GEN_608 : _GEN_2289; // @[Conditional.scala 40:58]
  wire [127:0] mask = _GEN_2298[127:0]; // @[dcache.scala 166:23]
  wire  _GEN_2504 = 4'h0 == blockIdx; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_326 = 2'h0 == _GEN_129 & 4'h0 == blockIdx | dirty_0_0; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_2507 = 4'h1 == blockIdx; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_327 = 2'h0 == _GEN_129 & 4'h1 == blockIdx | dirty_0_1; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_2510 = 4'h2 == blockIdx; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_328 = 2'h0 == _GEN_129 & 4'h2 == blockIdx | dirty_0_2; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_2513 = 4'h3 == blockIdx; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_329 = 2'h0 == _GEN_129 & 4'h3 == blockIdx | dirty_0_3; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_2516 = 4'h4 == blockIdx; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_330 = 2'h0 == _GEN_129 & 4'h4 == blockIdx | dirty_0_4; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_2519 = 4'h5 == blockIdx; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_331 = 2'h0 == _GEN_129 & 4'h5 == blockIdx | dirty_0_5; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_2522 = 4'h6 == blockIdx; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_332 = 2'h0 == _GEN_129 & 4'h6 == blockIdx | dirty_0_6; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_2525 = 4'h7 == blockIdx; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_333 = 2'h0 == _GEN_129 & 4'h7 == blockIdx | dirty_0_7; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_2528 = 4'h8 == blockIdx; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_334 = 2'h0 == _GEN_129 & 4'h8 == blockIdx | dirty_0_8; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_2531 = 4'h9 == blockIdx; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_335 = 2'h0 == _GEN_129 & 4'h9 == blockIdx | dirty_0_9; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_2534 = 4'ha == blockIdx; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_336 = 2'h0 == _GEN_129 & 4'ha == blockIdx | dirty_0_10; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_2537 = 4'hb == blockIdx; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_337 = 2'h0 == _GEN_129 & 4'hb == blockIdx | dirty_0_11; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_2540 = 4'hc == blockIdx; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_338 = 2'h0 == _GEN_129 & 4'hc == blockIdx | dirty_0_12; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_2543 = 4'hd == blockIdx; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_339 = 2'h0 == _GEN_129 & 4'hd == blockIdx | dirty_0_13; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_2546 = 4'he == blockIdx; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_340 = 2'h0 == _GEN_129 & 4'he == blockIdx | dirty_0_14; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_2549 = 4'hf == blockIdx; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_341 = 2'h0 == _GEN_129 & 4'hf == blockIdx | dirty_0_15; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_342 = 2'h1 == _GEN_129 & 4'h0 == blockIdx | dirty_1_0; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_343 = 2'h1 == _GEN_129 & 4'h1 == blockIdx | dirty_1_1; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_344 = 2'h1 == _GEN_129 & 4'h2 == blockIdx | dirty_1_2; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_345 = 2'h1 == _GEN_129 & 4'h3 == blockIdx | dirty_1_3; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_346 = 2'h1 == _GEN_129 & 4'h4 == blockIdx | dirty_1_4; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_347 = 2'h1 == _GEN_129 & 4'h5 == blockIdx | dirty_1_5; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_348 = 2'h1 == _GEN_129 & 4'h6 == blockIdx | dirty_1_6; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_349 = 2'h1 == _GEN_129 & 4'h7 == blockIdx | dirty_1_7; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_350 = 2'h1 == _GEN_129 & 4'h8 == blockIdx | dirty_1_8; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_351 = 2'h1 == _GEN_129 & 4'h9 == blockIdx | dirty_1_9; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_352 = 2'h1 == _GEN_129 & 4'ha == blockIdx | dirty_1_10; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_353 = 2'h1 == _GEN_129 & 4'hb == blockIdx | dirty_1_11; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_354 = 2'h1 == _GEN_129 & 4'hc == blockIdx | dirty_1_12; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_355 = 2'h1 == _GEN_129 & 4'hd == blockIdx | dirty_1_13; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_356 = 2'h1 == _GEN_129 & 4'he == blockIdx | dirty_1_14; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_357 = 2'h1 == _GEN_129 & 4'hf == blockIdx | dirty_1_15; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_358 = 2'h2 == _GEN_129 & 4'h0 == blockIdx | dirty_2_0; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_359 = 2'h2 == _GEN_129 & 4'h1 == blockIdx | dirty_2_1; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_360 = 2'h2 == _GEN_129 & 4'h2 == blockIdx | dirty_2_2; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_361 = 2'h2 == _GEN_129 & 4'h3 == blockIdx | dirty_2_3; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_362 = 2'h2 == _GEN_129 & 4'h4 == blockIdx | dirty_2_4; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_363 = 2'h2 == _GEN_129 & 4'h5 == blockIdx | dirty_2_5; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_364 = 2'h2 == _GEN_129 & 4'h6 == blockIdx | dirty_2_6; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_365 = 2'h2 == _GEN_129 & 4'h7 == blockIdx | dirty_2_7; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_366 = 2'h2 == _GEN_129 & 4'h8 == blockIdx | dirty_2_8; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_367 = 2'h2 == _GEN_129 & 4'h9 == blockIdx | dirty_2_9; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_368 = 2'h2 == _GEN_129 & 4'ha == blockIdx | dirty_2_10; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_369 = 2'h2 == _GEN_129 & 4'hb == blockIdx | dirty_2_11; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_370 = 2'h2 == _GEN_129 & 4'hc == blockIdx | dirty_2_12; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_371 = 2'h2 == _GEN_129 & 4'hd == blockIdx | dirty_2_13; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_372 = 2'h2 == _GEN_129 & 4'he == blockIdx | dirty_2_14; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_373 = 2'h2 == _GEN_129 & 4'hf == blockIdx | dirty_2_15; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_374 = 2'h3 == _GEN_129 & 4'h0 == blockIdx | dirty_3_0; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_375 = 2'h3 == _GEN_129 & 4'h1 == blockIdx | dirty_3_1; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_376 = 2'h3 == _GEN_129 & 4'h2 == blockIdx | dirty_3_2; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_377 = 2'h3 == _GEN_129 & 4'h3 == blockIdx | dirty_3_3; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_378 = 2'h3 == _GEN_129 & 4'h4 == blockIdx | dirty_3_4; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_379 = 2'h3 == _GEN_129 & 4'h5 == blockIdx | dirty_3_5; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_380 = 2'h3 == _GEN_129 & 4'h6 == blockIdx | dirty_3_6; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_381 = 2'h3 == _GEN_129 & 4'h7 == blockIdx | dirty_3_7; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_382 = 2'h3 == _GEN_129 & 4'h8 == blockIdx | dirty_3_8; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_383 = 2'h3 == _GEN_129 & 4'h9 == blockIdx | dirty_3_9; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_384 = 2'h3 == _GEN_129 & 4'ha == blockIdx | dirty_3_10; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_385 = 2'h3 == _GEN_129 & 4'hb == blockIdx | dirty_3_11; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_386 = 2'h3 == _GEN_129 & 4'hc == blockIdx | dirty_3_12; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_387 = 2'h3 == _GEN_129 & 4'hd == blockIdx | dirty_3_13; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_388 = 2'h3 == _GEN_129 & 4'he == blockIdx | dirty_3_14; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_389 = 2'h3 == _GEN_129 & 4'hf == blockIdx | dirty_3_15; // @[dcache.scala 214:34 dcache.scala 214:34 dcache.scala 94:26]
  wire  _GEN_390 = wen & _io_dc2sr0_addr_T_2 ? _GEN_326 : dirty_0_0; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_391 = wen & _io_dc2sr0_addr_T_2 ? _GEN_327 : dirty_0_1; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_392 = wen & _io_dc2sr0_addr_T_2 ? _GEN_328 : dirty_0_2; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_393 = wen & _io_dc2sr0_addr_T_2 ? _GEN_329 : dirty_0_3; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_394 = wen & _io_dc2sr0_addr_T_2 ? _GEN_330 : dirty_0_4; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_395 = wen & _io_dc2sr0_addr_T_2 ? _GEN_331 : dirty_0_5; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_396 = wen & _io_dc2sr0_addr_T_2 ? _GEN_332 : dirty_0_6; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_397 = wen & _io_dc2sr0_addr_T_2 ? _GEN_333 : dirty_0_7; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_398 = wen & _io_dc2sr0_addr_T_2 ? _GEN_334 : dirty_0_8; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_399 = wen & _io_dc2sr0_addr_T_2 ? _GEN_335 : dirty_0_9; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_400 = wen & _io_dc2sr0_addr_T_2 ? _GEN_336 : dirty_0_10; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_401 = wen & _io_dc2sr0_addr_T_2 ? _GEN_337 : dirty_0_11; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_402 = wen & _io_dc2sr0_addr_T_2 ? _GEN_338 : dirty_0_12; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_403 = wen & _io_dc2sr0_addr_T_2 ? _GEN_339 : dirty_0_13; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_404 = wen & _io_dc2sr0_addr_T_2 ? _GEN_340 : dirty_0_14; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_405 = wen & _io_dc2sr0_addr_T_2 ? _GEN_341 : dirty_0_15; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_406 = wen & _io_dc2sr0_addr_T_2 ? _GEN_342 : dirty_1_0; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_407 = wen & _io_dc2sr0_addr_T_2 ? _GEN_343 : dirty_1_1; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_408 = wen & _io_dc2sr0_addr_T_2 ? _GEN_344 : dirty_1_2; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_409 = wen & _io_dc2sr0_addr_T_2 ? _GEN_345 : dirty_1_3; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_410 = wen & _io_dc2sr0_addr_T_2 ? _GEN_346 : dirty_1_4; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_411 = wen & _io_dc2sr0_addr_T_2 ? _GEN_347 : dirty_1_5; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_412 = wen & _io_dc2sr0_addr_T_2 ? _GEN_348 : dirty_1_6; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_413 = wen & _io_dc2sr0_addr_T_2 ? _GEN_349 : dirty_1_7; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_414 = wen & _io_dc2sr0_addr_T_2 ? _GEN_350 : dirty_1_8; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_415 = wen & _io_dc2sr0_addr_T_2 ? _GEN_351 : dirty_1_9; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_416 = wen & _io_dc2sr0_addr_T_2 ? _GEN_352 : dirty_1_10; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_417 = wen & _io_dc2sr0_addr_T_2 ? _GEN_353 : dirty_1_11; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_418 = wen & _io_dc2sr0_addr_T_2 ? _GEN_354 : dirty_1_12; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_419 = wen & _io_dc2sr0_addr_T_2 ? _GEN_355 : dirty_1_13; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_420 = wen & _io_dc2sr0_addr_T_2 ? _GEN_356 : dirty_1_14; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_421 = wen & _io_dc2sr0_addr_T_2 ? _GEN_357 : dirty_1_15; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_422 = wen & _io_dc2sr0_addr_T_2 ? _GEN_358 : dirty_2_0; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_423 = wen & _io_dc2sr0_addr_T_2 ? _GEN_359 : dirty_2_1; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_424 = wen & _io_dc2sr0_addr_T_2 ? _GEN_360 : dirty_2_2; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_425 = wen & _io_dc2sr0_addr_T_2 ? _GEN_361 : dirty_2_3; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_426 = wen & _io_dc2sr0_addr_T_2 ? _GEN_362 : dirty_2_4; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_427 = wen & _io_dc2sr0_addr_T_2 ? _GEN_363 : dirty_2_5; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_428 = wen & _io_dc2sr0_addr_T_2 ? _GEN_364 : dirty_2_6; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_429 = wen & _io_dc2sr0_addr_T_2 ? _GEN_365 : dirty_2_7; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_430 = wen & _io_dc2sr0_addr_T_2 ? _GEN_366 : dirty_2_8; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_431 = wen & _io_dc2sr0_addr_T_2 ? _GEN_367 : dirty_2_9; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_432 = wen & _io_dc2sr0_addr_T_2 ? _GEN_368 : dirty_2_10; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_433 = wen & _io_dc2sr0_addr_T_2 ? _GEN_369 : dirty_2_11; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_434 = wen & _io_dc2sr0_addr_T_2 ? _GEN_370 : dirty_2_12; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_435 = wen & _io_dc2sr0_addr_T_2 ? _GEN_371 : dirty_2_13; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_436 = wen & _io_dc2sr0_addr_T_2 ? _GEN_372 : dirty_2_14; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_437 = wen & _io_dc2sr0_addr_T_2 ? _GEN_373 : dirty_2_15; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_438 = wen & _io_dc2sr0_addr_T_2 ? _GEN_374 : dirty_3_0; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_439 = wen & _io_dc2sr0_addr_T_2 ? _GEN_375 : dirty_3_1; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_440 = wen & _io_dc2sr0_addr_T_2 ? _GEN_376 : dirty_3_2; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_441 = wen & _io_dc2sr0_addr_T_2 ? _GEN_377 : dirty_3_3; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_442 = wen & _io_dc2sr0_addr_T_2 ? _GEN_378 : dirty_3_4; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_443 = wen & _io_dc2sr0_addr_T_2 ? _GEN_379 : dirty_3_5; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_444 = wen & _io_dc2sr0_addr_T_2 ? _GEN_380 : dirty_3_6; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_445 = wen & _io_dc2sr0_addr_T_2 ? _GEN_381 : dirty_3_7; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_446 = wen & _io_dc2sr0_addr_T_2 ? _GEN_382 : dirty_3_8; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_447 = wen & _io_dc2sr0_addr_T_2 ? _GEN_383 : dirty_3_9; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_448 = wen & _io_dc2sr0_addr_T_2 ? _GEN_384 : dirty_3_10; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_449 = wen & _io_dc2sr0_addr_T_2 ? _GEN_385 : dirty_3_11; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_450 = wen & _io_dc2sr0_addr_T_2 ? _GEN_386 : dirty_3_12; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_451 = wen & _io_dc2sr0_addr_T_2 ? _GEN_387 : dirty_3_13; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_452 = wen & _io_dc2sr0_addr_T_2 ? _GEN_388 : dirty_3_14; // @[dcache.scala 213:56 dcache.scala 94:26]
  wire  _GEN_453 = wen & _io_dc2sr0_addr_T_2 ? _GEN_389 : dirty_3_15; // @[dcache.scala 213:56 dcache.scala 94:26]
  reg  axiRaddrEn; // @[dcache.scala 218:34]
  reg  axiWaddrEn; // @[dcache.scala 221:34]
  wire  _GEN_2695 = 2'h0 == matchWay_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire  _GEN_2696 = 4'h1 == blockIdx_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_455 = 2'h0 == matchWay_r & 4'h1 == blockIdx_r ? tag_0_1 : tag_0_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire  _GEN_2698 = 4'h2 == blockIdx_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_456 = 2'h0 == matchWay_r & 4'h2 == blockIdx_r ? tag_0_2 : _GEN_455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire  _GEN_2700 = 4'h3 == blockIdx_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_457 = 2'h0 == matchWay_r & 4'h3 == blockIdx_r ? tag_0_3 : _GEN_456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire  _GEN_2702 = 4'h4 == blockIdx_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_458 = 2'h0 == matchWay_r & 4'h4 == blockIdx_r ? tag_0_4 : _GEN_457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire  _GEN_2704 = 4'h5 == blockIdx_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_459 = 2'h0 == matchWay_r & 4'h5 == blockIdx_r ? tag_0_5 : _GEN_458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire  _GEN_2706 = 4'h6 == blockIdx_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_460 = 2'h0 == matchWay_r & 4'h6 == blockIdx_r ? tag_0_6 : _GEN_459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire  _GEN_2708 = 4'h7 == blockIdx_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_461 = 2'h0 == matchWay_r & 4'h7 == blockIdx_r ? tag_0_7 : _GEN_460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire  _GEN_2710 = 4'h8 == blockIdx_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_462 = 2'h0 == matchWay_r & 4'h8 == blockIdx_r ? tag_0_8 : _GEN_461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire  _GEN_2712 = 4'h9 == blockIdx_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_463 = 2'h0 == matchWay_r & 4'h9 == blockIdx_r ? tag_0_9 : _GEN_462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire  _GEN_2714 = 4'ha == blockIdx_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_464 = 2'h0 == matchWay_r & 4'ha == blockIdx_r ? tag_0_10 : _GEN_463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire  _GEN_2716 = 4'hb == blockIdx_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_465 = 2'h0 == matchWay_r & 4'hb == blockIdx_r ? tag_0_11 : _GEN_464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire  _GEN_2718 = 4'hc == blockIdx_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_466 = 2'h0 == matchWay_r & 4'hc == blockIdx_r ? tag_0_12 : _GEN_465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire  _GEN_2720 = 4'hd == blockIdx_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_467 = 2'h0 == matchWay_r & 4'hd == blockIdx_r ? tag_0_13 : _GEN_466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire  _GEN_2722 = 4'he == blockIdx_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_468 = 2'h0 == matchWay_r & 4'he == blockIdx_r ? tag_0_14 : _GEN_467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire  _GEN_2724 = 4'hf == blockIdx_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_469 = 2'h0 == matchWay_r & 4'hf == blockIdx_r ? tag_0_15 : _GEN_468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire  _GEN_2726 = 4'h0 == blockIdx_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_470 = _rdata128_T & 4'h0 == blockIdx_r ? tag_1_0 : _GEN_469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_471 = _rdata128_T & 4'h1 == blockIdx_r ? tag_1_1 : _GEN_470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_472 = _rdata128_T & 4'h2 == blockIdx_r ? tag_1_2 : _GEN_471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_473 = _rdata128_T & 4'h3 == blockIdx_r ? tag_1_3 : _GEN_472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_474 = _rdata128_T & 4'h4 == blockIdx_r ? tag_1_4 : _GEN_473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_475 = _rdata128_T & 4'h5 == blockIdx_r ? tag_1_5 : _GEN_474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_476 = _rdata128_T & 4'h6 == blockIdx_r ? tag_1_6 : _GEN_475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_477 = _rdata128_T & 4'h7 == blockIdx_r ? tag_1_7 : _GEN_476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_478 = _rdata128_T & 4'h8 == blockIdx_r ? tag_1_8 : _GEN_477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_479 = _rdata128_T & 4'h9 == blockIdx_r ? tag_1_9 : _GEN_478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_480 = _rdata128_T & 4'ha == blockIdx_r ? tag_1_10 : _GEN_479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_481 = _rdata128_T & 4'hb == blockIdx_r ? tag_1_11 : _GEN_480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_482 = _rdata128_T & 4'hc == blockIdx_r ? tag_1_12 : _GEN_481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_483 = _rdata128_T & 4'hd == blockIdx_r ? tag_1_13 : _GEN_482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_484 = _rdata128_T & 4'he == blockIdx_r ? tag_1_14 : _GEN_483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_485 = _rdata128_T & 4'hf == blockIdx_r ? tag_1_15 : _GEN_484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_486 = _rdata128_T_2 & 4'h0 == blockIdx_r ? tag_2_0 : _GEN_485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_487 = _rdata128_T_2 & 4'h1 == blockIdx_r ? tag_2_1 : _GEN_486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_488 = _rdata128_T_2 & 4'h2 == blockIdx_r ? tag_2_2 : _GEN_487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_489 = _rdata128_T_2 & 4'h3 == blockIdx_r ? tag_2_3 : _GEN_488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_490 = _rdata128_T_2 & 4'h4 == blockIdx_r ? tag_2_4 : _GEN_489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_491 = _rdata128_T_2 & 4'h5 == blockIdx_r ? tag_2_5 : _GEN_490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_492 = _rdata128_T_2 & 4'h6 == blockIdx_r ? tag_2_6 : _GEN_491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_493 = _rdata128_T_2 & 4'h7 == blockIdx_r ? tag_2_7 : _GEN_492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_494 = _rdata128_T_2 & 4'h8 == blockIdx_r ? tag_2_8 : _GEN_493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_495 = _rdata128_T_2 & 4'h9 == blockIdx_r ? tag_2_9 : _GEN_494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_496 = _rdata128_T_2 & 4'ha == blockIdx_r ? tag_2_10 : _GEN_495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_497 = _rdata128_T_2 & 4'hb == blockIdx_r ? tag_2_11 : _GEN_496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_498 = _rdata128_T_2 & 4'hc == blockIdx_r ? tag_2_12 : _GEN_497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_499 = _rdata128_T_2 & 4'hd == blockIdx_r ? tag_2_13 : _GEN_498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_500 = _rdata128_T_2 & 4'he == blockIdx_r ? tag_2_14 : _GEN_499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_501 = _rdata128_T_2 & 4'hf == blockIdx_r ? tag_2_15 : _GEN_500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_502 = _rdata128_T_4 & 4'h0 == blockIdx_r ? tag_3_0 : _GEN_501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_503 = _rdata128_T_4 & 4'h1 == blockIdx_r ? tag_3_1 : _GEN_502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_504 = _rdata128_T_4 & 4'h2 == blockIdx_r ? tag_3_2 : _GEN_503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_505 = _rdata128_T_4 & 4'h3 == blockIdx_r ? tag_3_3 : _GEN_504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_506 = _rdata128_T_4 & 4'h4 == blockIdx_r ? tag_3_4 : _GEN_505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_507 = _rdata128_T_4 & 4'h5 == blockIdx_r ? tag_3_5 : _GEN_506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_508 = _rdata128_T_4 & 4'h6 == blockIdx_r ? tag_3_6 : _GEN_507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_509 = _rdata128_T_4 & 4'h7 == blockIdx_r ? tag_3_7 : _GEN_508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_510 = _rdata128_T_4 & 4'h8 == blockIdx_r ? tag_3_8 : _GEN_509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_511 = _rdata128_T_4 & 4'h9 == blockIdx_r ? tag_3_9 : _GEN_510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_512 = _rdata128_T_4 & 4'ha == blockIdx_r ? tag_3_10 : _GEN_511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_513 = _rdata128_T_4 & 4'hb == blockIdx_r ? tag_3_11 : _GEN_512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_514 = _rdata128_T_4 & 4'hc == blockIdx_r ? tag_3_12 : _GEN_513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_515 = _rdata128_T_4 & 4'hd == blockIdx_r ? tag_3_13 : _GEN_514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_516 = _rdata128_T_4 & 4'he == blockIdx_r ? tag_3_14 : _GEN_515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_517 = _rdata128_T_4 & 4'hf == blockIdx_r ? tag_3_15 : _GEN_516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [25:0] axiWaddr_hi = {_GEN_517,blockIdx_r}; // @[Cat.scala 30:58]
  reg  axiWdataEn; // @[dcache.scala 224:34]
  wire [2:0] _GEN_518 = cur_mode_sl == 2'h3 ? 3'h5 : state; // @[dcache.scala 234:42 dcache.scala 235:27 dcache.scala 153:24]
  wire  _GEN_524 = 2'h0 == matchWay & _GEN_2507 ? dirty_0_1 : dirty_0_0; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_525 = 2'h0 == matchWay & _GEN_2510 ? dirty_0_2 : _GEN_524; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_526 = 2'h0 == matchWay & _GEN_2513 ? dirty_0_3 : _GEN_525; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_527 = 2'h0 == matchWay & _GEN_2516 ? dirty_0_4 : _GEN_526; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_528 = 2'h0 == matchWay & _GEN_2519 ? dirty_0_5 : _GEN_527; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_529 = 2'h0 == matchWay & _GEN_2522 ? dirty_0_6 : _GEN_528; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_530 = 2'h0 == matchWay & _GEN_2525 ? dirty_0_7 : _GEN_529; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_531 = 2'h0 == matchWay & _GEN_2528 ? dirty_0_8 : _GEN_530; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_532 = 2'h0 == matchWay & _GEN_2531 ? dirty_0_9 : _GEN_531; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_533 = 2'h0 == matchWay & _GEN_2534 ? dirty_0_10 : _GEN_532; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_534 = 2'h0 == matchWay & _GEN_2537 ? dirty_0_11 : _GEN_533; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_535 = 2'h0 == matchWay & _GEN_2540 ? dirty_0_12 : _GEN_534; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_536 = 2'h0 == matchWay & _GEN_2543 ? dirty_0_13 : _GEN_535; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_537 = 2'h0 == matchWay & _GEN_2546 ? dirty_0_14 : _GEN_536; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_538 = 2'h0 == matchWay & _GEN_2549 ? dirty_0_15 : _GEN_537; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_539 = 2'h1 == matchWay & _GEN_2504 ? dirty_1_0 : _GEN_538; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_540 = 2'h1 == matchWay & _GEN_2507 ? dirty_1_1 : _GEN_539; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_541 = 2'h1 == matchWay & _GEN_2510 ? dirty_1_2 : _GEN_540; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_542 = 2'h1 == matchWay & _GEN_2513 ? dirty_1_3 : _GEN_541; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_543 = 2'h1 == matchWay & _GEN_2516 ? dirty_1_4 : _GEN_542; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_544 = 2'h1 == matchWay & _GEN_2519 ? dirty_1_5 : _GEN_543; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_545 = 2'h1 == matchWay & _GEN_2522 ? dirty_1_6 : _GEN_544; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_546 = 2'h1 == matchWay & _GEN_2525 ? dirty_1_7 : _GEN_545; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_547 = 2'h1 == matchWay & _GEN_2528 ? dirty_1_8 : _GEN_546; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_548 = 2'h1 == matchWay & _GEN_2531 ? dirty_1_9 : _GEN_547; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_549 = 2'h1 == matchWay & _GEN_2534 ? dirty_1_10 : _GEN_548; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_550 = 2'h1 == matchWay & _GEN_2537 ? dirty_1_11 : _GEN_549; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_551 = 2'h1 == matchWay & _GEN_2540 ? dirty_1_12 : _GEN_550; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_552 = 2'h1 == matchWay & _GEN_2543 ? dirty_1_13 : _GEN_551; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_553 = 2'h1 == matchWay & _GEN_2546 ? dirty_1_14 : _GEN_552; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_554 = 2'h1 == matchWay & _GEN_2549 ? dirty_1_15 : _GEN_553; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_555 = 2'h2 == matchWay & _GEN_2504 ? dirty_2_0 : _GEN_554; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_556 = 2'h2 == matchWay & _GEN_2507 ? dirty_2_1 : _GEN_555; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_557 = 2'h2 == matchWay & _GEN_2510 ? dirty_2_2 : _GEN_556; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_558 = 2'h2 == matchWay & _GEN_2513 ? dirty_2_3 : _GEN_557; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_559 = 2'h2 == matchWay & _GEN_2516 ? dirty_2_4 : _GEN_558; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_560 = 2'h2 == matchWay & _GEN_2519 ? dirty_2_5 : _GEN_559; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_561 = 2'h2 == matchWay & _GEN_2522 ? dirty_2_6 : _GEN_560; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_562 = 2'h2 == matchWay & _GEN_2525 ? dirty_2_7 : _GEN_561; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_563 = 2'h2 == matchWay & _GEN_2528 ? dirty_2_8 : _GEN_562; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_564 = 2'h2 == matchWay & _GEN_2531 ? dirty_2_9 : _GEN_563; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_565 = 2'h2 == matchWay & _GEN_2534 ? dirty_2_10 : _GEN_564; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_566 = 2'h2 == matchWay & _GEN_2537 ? dirty_2_11 : _GEN_565; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_567 = 2'h2 == matchWay & _GEN_2540 ? dirty_2_12 : _GEN_566; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_568 = 2'h2 == matchWay & _GEN_2543 ? dirty_2_13 : _GEN_567; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_569 = 2'h2 == matchWay & _GEN_2546 ? dirty_2_14 : _GEN_568; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_570 = 2'h2 == matchWay & _GEN_2549 ? dirty_2_15 : _GEN_569; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_571 = 2'h3 == matchWay & _GEN_2504 ? dirty_3_0 : _GEN_570; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_572 = 2'h3 == matchWay & _GEN_2507 ? dirty_3_1 : _GEN_571; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_573 = 2'h3 == matchWay & _GEN_2510 ? dirty_3_2 : _GEN_572; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_574 = 2'h3 == matchWay & _GEN_2513 ? dirty_3_3 : _GEN_573; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_575 = 2'h3 == matchWay & _GEN_2516 ? dirty_3_4 : _GEN_574; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_576 = 2'h3 == matchWay & _GEN_2519 ? dirty_3_5 : _GEN_575; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_577 = 2'h3 == matchWay & _GEN_2522 ? dirty_3_6 : _GEN_576; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_578 = 2'h3 == matchWay & _GEN_2525 ? dirty_3_7 : _GEN_577; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_579 = 2'h3 == matchWay & _GEN_2528 ? dirty_3_8 : _GEN_578; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_580 = 2'h3 == matchWay & _GEN_2531 ? dirty_3_9 : _GEN_579; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_581 = 2'h3 == matchWay & _GEN_2534 ? dirty_3_10 : _GEN_580; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_582 = 2'h3 == matchWay & _GEN_2537 ? dirty_3_11 : _GEN_581; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_583 = 2'h3 == matchWay & _GEN_2540 ? dirty_3_12 : _GEN_582; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_584 = 2'h3 == matchWay & _GEN_2543 ? dirty_3_13 : _GEN_583; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_585 = 2'h3 == matchWay & _GEN_2546 ? dirty_3_14 : _GEN_584; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire  _GEN_586 = 2'h3 == matchWay & _GEN_2549 ? dirty_3_15 : _GEN_585; // @[dcache.scala 245:31 dcache.scala 245:31]
  wire [2:0] _GEN_587 = _GEN_586 ? 3'h3 : 3'h1; // @[dcache.scala 245:31 dcache.scala 246:27 dcache.scala 249:27]
  wire  _GEN_588 = _GEN_586 | axiWaddrEn; // @[dcache.scala 245:31 dcache.scala 247:32 dcache.scala 221:34]
  wire  _GEN_589 = _GEN_586 ? axiRaddrEn : 1'h1; // @[dcache.scala 245:31 dcache.scala 218:34 dcache.scala 250:32]
  wire [2:0] _GEN_590 = cacheHit ? _GEN_518 : _GEN_587; // @[dcache.scala 233:33]
  wire  _GEN_592 = cacheHit ? _T_73 : 1'h1; // @[dcache.scala 233:33 dcache.scala 253:25]
  wire  _GEN_595 = cacheHit ? axiWaddrEn : _GEN_588; // @[dcache.scala 233:33 dcache.scala 221:34]
  wire  _GEN_596 = cacheHit ? axiRaddrEn : _GEN_589; // @[dcache.scala 233:33 dcache.scala 218:34]
  wire  _GEN_598 = ~hs_in & _io_dcRW_ready_T ? 1'h0 : cacheHit; // @[dcache.scala 231:42 dcache.scala 102:13]
  wire  _GEN_605 = flush_r | io_flush ? 1'h0 : _GEN_598; // @[dcache.scala 229:38 dcache.scala 102:13]
  wire  _GEN_613 = axiRaddrEn & io_dataAxi_ra_ready | axiRdataEn; // @[dcache.scala 258:52 dcache.scala 261:28 dcache.scala 220:34]
  wire [2:0] _offset_T_1 = offset + 3'h1; // @[dcache.scala 266:34]
  wire [63:0] _GEN_615 = offset[0] ? rdatabuf : io_dataAxi_rd_bits_data; // @[dcache.scala 267:32 dcache.scala 112:34 dcache.scala 270:30]
  wire  _GEN_2948 = 4'h0 == pre_blockIdx; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_616 = _GEN_2695 & 4'h0 == pre_blockIdx ? pre_tag : tag_0_0; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire  _GEN_2950 = 4'h1 == pre_blockIdx; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_617 = _GEN_2695 & 4'h1 == pre_blockIdx ? pre_tag : tag_0_1; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire  _GEN_2952 = 4'h2 == pre_blockIdx; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_618 = _GEN_2695 & 4'h2 == pre_blockIdx ? pre_tag : tag_0_2; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire  _GEN_2954 = 4'h3 == pre_blockIdx; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_619 = _GEN_2695 & 4'h3 == pre_blockIdx ? pre_tag : tag_0_3; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire  _GEN_2956 = 4'h4 == pre_blockIdx; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_620 = _GEN_2695 & 4'h4 == pre_blockIdx ? pre_tag : tag_0_4; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire  _GEN_2958 = 4'h5 == pre_blockIdx; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_621 = _GEN_2695 & 4'h5 == pre_blockIdx ? pre_tag : tag_0_5; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire  _GEN_2960 = 4'h6 == pre_blockIdx; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_622 = _GEN_2695 & 4'h6 == pre_blockIdx ? pre_tag : tag_0_6; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire  _GEN_2962 = 4'h7 == pre_blockIdx; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_623 = _GEN_2695 & 4'h7 == pre_blockIdx ? pre_tag : tag_0_7; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire  _GEN_2964 = 4'h8 == pre_blockIdx; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_624 = _GEN_2695 & 4'h8 == pre_blockIdx ? pre_tag : tag_0_8; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire  _GEN_2966 = 4'h9 == pre_blockIdx; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_625 = _GEN_2695 & 4'h9 == pre_blockIdx ? pre_tag : tag_0_9; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire  _GEN_2968 = 4'ha == pre_blockIdx; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_626 = _GEN_2695 & 4'ha == pre_blockIdx ? pre_tag : tag_0_10; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire  _GEN_2970 = 4'hb == pre_blockIdx; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_627 = _GEN_2695 & 4'hb == pre_blockIdx ? pre_tag : tag_0_11; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire  _GEN_2972 = 4'hc == pre_blockIdx; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_628 = _GEN_2695 & 4'hc == pre_blockIdx ? pre_tag : tag_0_12; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire  _GEN_2974 = 4'hd == pre_blockIdx; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_629 = _GEN_2695 & 4'hd == pre_blockIdx ? pre_tag : tag_0_13; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire  _GEN_2976 = 4'he == pre_blockIdx; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_630 = _GEN_2695 & 4'he == pre_blockIdx ? pre_tag : tag_0_14; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire  _GEN_2978 = 4'hf == pre_blockIdx; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_631 = _GEN_2695 & 4'hf == pre_blockIdx ? pre_tag : tag_0_15; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_632 = _rdata128_T & 4'h0 == pre_blockIdx ? pre_tag : tag_1_0; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_633 = _rdata128_T & 4'h1 == pre_blockIdx ? pre_tag : tag_1_1; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_634 = _rdata128_T & 4'h2 == pre_blockIdx ? pre_tag : tag_1_2; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_635 = _rdata128_T & 4'h3 == pre_blockIdx ? pre_tag : tag_1_3; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_636 = _rdata128_T & 4'h4 == pre_blockIdx ? pre_tag : tag_1_4; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_637 = _rdata128_T & 4'h5 == pre_blockIdx ? pre_tag : tag_1_5; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_638 = _rdata128_T & 4'h6 == pre_blockIdx ? pre_tag : tag_1_6; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_639 = _rdata128_T & 4'h7 == pre_blockIdx ? pre_tag : tag_1_7; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_640 = _rdata128_T & 4'h8 == pre_blockIdx ? pre_tag : tag_1_8; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_641 = _rdata128_T & 4'h9 == pre_blockIdx ? pre_tag : tag_1_9; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_642 = _rdata128_T & 4'ha == pre_blockIdx ? pre_tag : tag_1_10; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_643 = _rdata128_T & 4'hb == pre_blockIdx ? pre_tag : tag_1_11; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_644 = _rdata128_T & 4'hc == pre_blockIdx ? pre_tag : tag_1_12; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_645 = _rdata128_T & 4'hd == pre_blockIdx ? pre_tag : tag_1_13; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_646 = _rdata128_T & 4'he == pre_blockIdx ? pre_tag : tag_1_14; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_647 = _rdata128_T & 4'hf == pre_blockIdx ? pre_tag : tag_1_15; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_648 = _rdata128_T_2 & 4'h0 == pre_blockIdx ? pre_tag : tag_2_0; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_649 = _rdata128_T_2 & 4'h1 == pre_blockIdx ? pre_tag : tag_2_1; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_650 = _rdata128_T_2 & 4'h2 == pre_blockIdx ? pre_tag : tag_2_2; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_651 = _rdata128_T_2 & 4'h3 == pre_blockIdx ? pre_tag : tag_2_3; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_652 = _rdata128_T_2 & 4'h4 == pre_blockIdx ? pre_tag : tag_2_4; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_653 = _rdata128_T_2 & 4'h5 == pre_blockIdx ? pre_tag : tag_2_5; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_654 = _rdata128_T_2 & 4'h6 == pre_blockIdx ? pre_tag : tag_2_6; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_655 = _rdata128_T_2 & 4'h7 == pre_blockIdx ? pre_tag : tag_2_7; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_656 = _rdata128_T_2 & 4'h8 == pre_blockIdx ? pre_tag : tag_2_8; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_657 = _rdata128_T_2 & 4'h9 == pre_blockIdx ? pre_tag : tag_2_9; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_658 = _rdata128_T_2 & 4'ha == pre_blockIdx ? pre_tag : tag_2_10; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_659 = _rdata128_T_2 & 4'hb == pre_blockIdx ? pre_tag : tag_2_11; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_660 = _rdata128_T_2 & 4'hc == pre_blockIdx ? pre_tag : tag_2_12; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_661 = _rdata128_T_2 & 4'hd == pre_blockIdx ? pre_tag : tag_2_13; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_662 = _rdata128_T_2 & 4'he == pre_blockIdx ? pre_tag : tag_2_14; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_663 = _rdata128_T_2 & 4'hf == pre_blockIdx ? pre_tag : tag_2_15; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_664 = _rdata128_T_4 & 4'h0 == pre_blockIdx ? pre_tag : tag_3_0; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_665 = _rdata128_T_4 & 4'h1 == pre_blockIdx ? pre_tag : tag_3_1; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_666 = _rdata128_T_4 & 4'h2 == pre_blockIdx ? pre_tag : tag_3_2; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_667 = _rdata128_T_4 & 4'h3 == pre_blockIdx ? pre_tag : tag_3_3; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_668 = _rdata128_T_4 & 4'h4 == pre_blockIdx ? pre_tag : tag_3_4; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_669 = _rdata128_T_4 & 4'h5 == pre_blockIdx ? pre_tag : tag_3_5; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_670 = _rdata128_T_4 & 4'h6 == pre_blockIdx ? pre_tag : tag_3_6; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_671 = _rdata128_T_4 & 4'h7 == pre_blockIdx ? pre_tag : tag_3_7; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_672 = _rdata128_T_4 & 4'h8 == pre_blockIdx ? pre_tag : tag_3_8; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_673 = _rdata128_T_4 & 4'h9 == pre_blockIdx ? pre_tag : tag_3_9; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_674 = _rdata128_T_4 & 4'ha == pre_blockIdx ? pre_tag : tag_3_10; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_675 = _rdata128_T_4 & 4'hb == pre_blockIdx ? pre_tag : tag_3_11; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_676 = _rdata128_T_4 & 4'hc == pre_blockIdx ? pre_tag : tag_3_12; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_677 = _rdata128_T_4 & 4'hd == pre_blockIdx ? pre_tag : tag_3_13; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_678 = _rdata128_T_4 & 4'he == pre_blockIdx ? pre_tag : tag_3_14; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire [21:0] _GEN_679 = _rdata128_T_4 & 4'hf == pre_blockIdx ? pre_tag : tag_3_15; // @[dcache.scala 274:51 dcache.scala 274:51 dcache.scala 92:26]
  wire  _GEN_680 = _GEN_2695 & _GEN_2948 | valid_0_0; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_681 = _GEN_2695 & _GEN_2950 | valid_0_1; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_682 = _GEN_2695 & _GEN_2952 | valid_0_2; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_683 = _GEN_2695 & _GEN_2954 | valid_0_3; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_684 = _GEN_2695 & _GEN_2956 | valid_0_4; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_685 = _GEN_2695 & _GEN_2958 | valid_0_5; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_686 = _GEN_2695 & _GEN_2960 | valid_0_6; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_687 = _GEN_2695 & _GEN_2962 | valid_0_7; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_688 = _GEN_2695 & _GEN_2964 | valid_0_8; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_689 = _GEN_2695 & _GEN_2966 | valid_0_9; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_690 = _GEN_2695 & _GEN_2968 | valid_0_10; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_691 = _GEN_2695 & _GEN_2970 | valid_0_11; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_692 = _GEN_2695 & _GEN_2972 | valid_0_12; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_693 = _GEN_2695 & _GEN_2974 | valid_0_13; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_694 = _GEN_2695 & _GEN_2976 | valid_0_14; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_695 = _GEN_2695 & _GEN_2978 | valid_0_15; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_696 = _rdata128_T & _GEN_2948 | valid_1_0; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_697 = _rdata128_T & _GEN_2950 | valid_1_1; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_698 = _rdata128_T & _GEN_2952 | valid_1_2; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_699 = _rdata128_T & _GEN_2954 | valid_1_3; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_700 = _rdata128_T & _GEN_2956 | valid_1_4; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_701 = _rdata128_T & _GEN_2958 | valid_1_5; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_702 = _rdata128_T & _GEN_2960 | valid_1_6; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_703 = _rdata128_T & _GEN_2962 | valid_1_7; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_704 = _rdata128_T & _GEN_2964 | valid_1_8; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_705 = _rdata128_T & _GEN_2966 | valid_1_9; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_706 = _rdata128_T & _GEN_2968 | valid_1_10; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_707 = _rdata128_T & _GEN_2970 | valid_1_11; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_708 = _rdata128_T & _GEN_2972 | valid_1_12; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_709 = _rdata128_T & _GEN_2974 | valid_1_13; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_710 = _rdata128_T & _GEN_2976 | valid_1_14; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_711 = _rdata128_T & _GEN_2978 | valid_1_15; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_712 = _rdata128_T_2 & _GEN_2948 | valid_2_0; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_713 = _rdata128_T_2 & _GEN_2950 | valid_2_1; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_714 = _rdata128_T_2 & _GEN_2952 | valid_2_2; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_715 = _rdata128_T_2 & _GEN_2954 | valid_2_3; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_716 = _rdata128_T_2 & _GEN_2956 | valid_2_4; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_717 = _rdata128_T_2 & _GEN_2958 | valid_2_5; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_718 = _rdata128_T_2 & _GEN_2960 | valid_2_6; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_719 = _rdata128_T_2 & _GEN_2962 | valid_2_7; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_720 = _rdata128_T_2 & _GEN_2964 | valid_2_8; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_721 = _rdata128_T_2 & _GEN_2966 | valid_2_9; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_722 = _rdata128_T_2 & _GEN_2968 | valid_2_10; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_723 = _rdata128_T_2 & _GEN_2970 | valid_2_11; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_724 = _rdata128_T_2 & _GEN_2972 | valid_2_12; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_725 = _rdata128_T_2 & _GEN_2974 | valid_2_13; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_726 = _rdata128_T_2 & _GEN_2976 | valid_2_14; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_727 = _rdata128_T_2 & _GEN_2978 | valid_2_15; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_728 = _rdata128_T_4 & _GEN_2948 | valid_3_0; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_729 = _rdata128_T_4 & _GEN_2950 | valid_3_1; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_730 = _rdata128_T_4 & _GEN_2952 | valid_3_2; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_731 = _rdata128_T_4 & _GEN_2954 | valid_3_3; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_732 = _rdata128_T_4 & _GEN_2956 | valid_3_4; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_733 = _rdata128_T_4 & _GEN_2958 | valid_3_5; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_734 = _rdata128_T_4 & _GEN_2960 | valid_3_6; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_735 = _rdata128_T_4 & _GEN_2962 | valid_3_7; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_736 = _rdata128_T_4 & _GEN_2964 | valid_3_8; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_737 = _rdata128_T_4 & _GEN_2966 | valid_3_9; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_738 = _rdata128_T_4 & _GEN_2968 | valid_3_10; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_739 = _rdata128_T_4 & _GEN_2970 | valid_3_11; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_740 = _rdata128_T_4 & _GEN_2972 | valid_3_12; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_741 = _rdata128_T_4 & _GEN_2974 | valid_3_13; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_742 = _rdata128_T_4 & _GEN_2976 | valid_3_14; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_743 = _rdata128_T_4 & _GEN_2978 | valid_3_15; // @[dcache.scala 275:53 dcache.scala 275:53 dcache.scala 93:26]
  wire  _GEN_744 = io_dataAxi_rd_bits_last ? 1'h0 : axiRdataEn; // @[dcache.scala 272:46 dcache.scala 273:32 dcache.scala 220:34]
  wire [21:0] _GEN_745 = io_dataAxi_rd_bits_last ? _GEN_616 : tag_0_0; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_746 = io_dataAxi_rd_bits_last ? _GEN_617 : tag_0_1; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_747 = io_dataAxi_rd_bits_last ? _GEN_618 : tag_0_2; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_748 = io_dataAxi_rd_bits_last ? _GEN_619 : tag_0_3; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_749 = io_dataAxi_rd_bits_last ? _GEN_620 : tag_0_4; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_750 = io_dataAxi_rd_bits_last ? _GEN_621 : tag_0_5; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_751 = io_dataAxi_rd_bits_last ? _GEN_622 : tag_0_6; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_752 = io_dataAxi_rd_bits_last ? _GEN_623 : tag_0_7; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_753 = io_dataAxi_rd_bits_last ? _GEN_624 : tag_0_8; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_754 = io_dataAxi_rd_bits_last ? _GEN_625 : tag_0_9; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_755 = io_dataAxi_rd_bits_last ? _GEN_626 : tag_0_10; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_756 = io_dataAxi_rd_bits_last ? _GEN_627 : tag_0_11; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_757 = io_dataAxi_rd_bits_last ? _GEN_628 : tag_0_12; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_758 = io_dataAxi_rd_bits_last ? _GEN_629 : tag_0_13; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_759 = io_dataAxi_rd_bits_last ? _GEN_630 : tag_0_14; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_760 = io_dataAxi_rd_bits_last ? _GEN_631 : tag_0_15; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_761 = io_dataAxi_rd_bits_last ? _GEN_632 : tag_1_0; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_762 = io_dataAxi_rd_bits_last ? _GEN_633 : tag_1_1; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_763 = io_dataAxi_rd_bits_last ? _GEN_634 : tag_1_2; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_764 = io_dataAxi_rd_bits_last ? _GEN_635 : tag_1_3; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_765 = io_dataAxi_rd_bits_last ? _GEN_636 : tag_1_4; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_766 = io_dataAxi_rd_bits_last ? _GEN_637 : tag_1_5; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_767 = io_dataAxi_rd_bits_last ? _GEN_638 : tag_1_6; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_768 = io_dataAxi_rd_bits_last ? _GEN_639 : tag_1_7; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_769 = io_dataAxi_rd_bits_last ? _GEN_640 : tag_1_8; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_770 = io_dataAxi_rd_bits_last ? _GEN_641 : tag_1_9; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_771 = io_dataAxi_rd_bits_last ? _GEN_642 : tag_1_10; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_772 = io_dataAxi_rd_bits_last ? _GEN_643 : tag_1_11; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_773 = io_dataAxi_rd_bits_last ? _GEN_644 : tag_1_12; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_774 = io_dataAxi_rd_bits_last ? _GEN_645 : tag_1_13; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_775 = io_dataAxi_rd_bits_last ? _GEN_646 : tag_1_14; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_776 = io_dataAxi_rd_bits_last ? _GEN_647 : tag_1_15; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_777 = io_dataAxi_rd_bits_last ? _GEN_648 : tag_2_0; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_778 = io_dataAxi_rd_bits_last ? _GEN_649 : tag_2_1; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_779 = io_dataAxi_rd_bits_last ? _GEN_650 : tag_2_2; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_780 = io_dataAxi_rd_bits_last ? _GEN_651 : tag_2_3; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_781 = io_dataAxi_rd_bits_last ? _GEN_652 : tag_2_4; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_782 = io_dataAxi_rd_bits_last ? _GEN_653 : tag_2_5; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_783 = io_dataAxi_rd_bits_last ? _GEN_654 : tag_2_6; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_784 = io_dataAxi_rd_bits_last ? _GEN_655 : tag_2_7; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_785 = io_dataAxi_rd_bits_last ? _GEN_656 : tag_2_8; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_786 = io_dataAxi_rd_bits_last ? _GEN_657 : tag_2_9; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_787 = io_dataAxi_rd_bits_last ? _GEN_658 : tag_2_10; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_788 = io_dataAxi_rd_bits_last ? _GEN_659 : tag_2_11; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_789 = io_dataAxi_rd_bits_last ? _GEN_660 : tag_2_12; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_790 = io_dataAxi_rd_bits_last ? _GEN_661 : tag_2_13; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_791 = io_dataAxi_rd_bits_last ? _GEN_662 : tag_2_14; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_792 = io_dataAxi_rd_bits_last ? _GEN_663 : tag_2_15; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_793 = io_dataAxi_rd_bits_last ? _GEN_664 : tag_3_0; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_794 = io_dataAxi_rd_bits_last ? _GEN_665 : tag_3_1; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_795 = io_dataAxi_rd_bits_last ? _GEN_666 : tag_3_2; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_796 = io_dataAxi_rd_bits_last ? _GEN_667 : tag_3_3; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_797 = io_dataAxi_rd_bits_last ? _GEN_668 : tag_3_4; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_798 = io_dataAxi_rd_bits_last ? _GEN_669 : tag_3_5; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_799 = io_dataAxi_rd_bits_last ? _GEN_670 : tag_3_6; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_800 = io_dataAxi_rd_bits_last ? _GEN_671 : tag_3_7; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_801 = io_dataAxi_rd_bits_last ? _GEN_672 : tag_3_8; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_802 = io_dataAxi_rd_bits_last ? _GEN_673 : tag_3_9; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_803 = io_dataAxi_rd_bits_last ? _GEN_674 : tag_3_10; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_804 = io_dataAxi_rd_bits_last ? _GEN_675 : tag_3_11; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_805 = io_dataAxi_rd_bits_last ? _GEN_676 : tag_3_12; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_806 = io_dataAxi_rd_bits_last ? _GEN_677 : tag_3_13; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_807 = io_dataAxi_rd_bits_last ? _GEN_678 : tag_3_14; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire [21:0] _GEN_808 = io_dataAxi_rd_bits_last ? _GEN_679 : tag_3_15; // @[dcache.scala 272:46 dcache.scala 92:26]
  wire  _GEN_809 = io_dataAxi_rd_bits_last ? _GEN_680 : valid_0_0; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_810 = io_dataAxi_rd_bits_last ? _GEN_681 : valid_0_1; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_811 = io_dataAxi_rd_bits_last ? _GEN_682 : valid_0_2; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_812 = io_dataAxi_rd_bits_last ? _GEN_683 : valid_0_3; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_813 = io_dataAxi_rd_bits_last ? _GEN_684 : valid_0_4; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_814 = io_dataAxi_rd_bits_last ? _GEN_685 : valid_0_5; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_815 = io_dataAxi_rd_bits_last ? _GEN_686 : valid_0_6; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_816 = io_dataAxi_rd_bits_last ? _GEN_687 : valid_0_7; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_817 = io_dataAxi_rd_bits_last ? _GEN_688 : valid_0_8; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_818 = io_dataAxi_rd_bits_last ? _GEN_689 : valid_0_9; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_819 = io_dataAxi_rd_bits_last ? _GEN_690 : valid_0_10; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_820 = io_dataAxi_rd_bits_last ? _GEN_691 : valid_0_11; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_821 = io_dataAxi_rd_bits_last ? _GEN_692 : valid_0_12; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_822 = io_dataAxi_rd_bits_last ? _GEN_693 : valid_0_13; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_823 = io_dataAxi_rd_bits_last ? _GEN_694 : valid_0_14; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_824 = io_dataAxi_rd_bits_last ? _GEN_695 : valid_0_15; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_825 = io_dataAxi_rd_bits_last ? _GEN_696 : valid_1_0; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_826 = io_dataAxi_rd_bits_last ? _GEN_697 : valid_1_1; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_827 = io_dataAxi_rd_bits_last ? _GEN_698 : valid_1_2; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_828 = io_dataAxi_rd_bits_last ? _GEN_699 : valid_1_3; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_829 = io_dataAxi_rd_bits_last ? _GEN_700 : valid_1_4; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_830 = io_dataAxi_rd_bits_last ? _GEN_701 : valid_1_5; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_831 = io_dataAxi_rd_bits_last ? _GEN_702 : valid_1_6; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_832 = io_dataAxi_rd_bits_last ? _GEN_703 : valid_1_7; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_833 = io_dataAxi_rd_bits_last ? _GEN_704 : valid_1_8; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_834 = io_dataAxi_rd_bits_last ? _GEN_705 : valid_1_9; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_835 = io_dataAxi_rd_bits_last ? _GEN_706 : valid_1_10; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_836 = io_dataAxi_rd_bits_last ? _GEN_707 : valid_1_11; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_837 = io_dataAxi_rd_bits_last ? _GEN_708 : valid_1_12; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_838 = io_dataAxi_rd_bits_last ? _GEN_709 : valid_1_13; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_839 = io_dataAxi_rd_bits_last ? _GEN_710 : valid_1_14; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_840 = io_dataAxi_rd_bits_last ? _GEN_711 : valid_1_15; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_841 = io_dataAxi_rd_bits_last ? _GEN_712 : valid_2_0; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_842 = io_dataAxi_rd_bits_last ? _GEN_713 : valid_2_1; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_843 = io_dataAxi_rd_bits_last ? _GEN_714 : valid_2_2; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_844 = io_dataAxi_rd_bits_last ? _GEN_715 : valid_2_3; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_845 = io_dataAxi_rd_bits_last ? _GEN_716 : valid_2_4; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_846 = io_dataAxi_rd_bits_last ? _GEN_717 : valid_2_5; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_847 = io_dataAxi_rd_bits_last ? _GEN_718 : valid_2_6; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_848 = io_dataAxi_rd_bits_last ? _GEN_719 : valid_2_7; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_849 = io_dataAxi_rd_bits_last ? _GEN_720 : valid_2_8; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_850 = io_dataAxi_rd_bits_last ? _GEN_721 : valid_2_9; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_851 = io_dataAxi_rd_bits_last ? _GEN_722 : valid_2_10; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_852 = io_dataAxi_rd_bits_last ? _GEN_723 : valid_2_11; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_853 = io_dataAxi_rd_bits_last ? _GEN_724 : valid_2_12; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_854 = io_dataAxi_rd_bits_last ? _GEN_725 : valid_2_13; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_855 = io_dataAxi_rd_bits_last ? _GEN_726 : valid_2_14; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_856 = io_dataAxi_rd_bits_last ? _GEN_727 : valid_2_15; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_857 = io_dataAxi_rd_bits_last ? _GEN_728 : valid_3_0; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_858 = io_dataAxi_rd_bits_last ? _GEN_729 : valid_3_1; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_859 = io_dataAxi_rd_bits_last ? _GEN_730 : valid_3_2; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_860 = io_dataAxi_rd_bits_last ? _GEN_731 : valid_3_3; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_861 = io_dataAxi_rd_bits_last ? _GEN_732 : valid_3_4; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_862 = io_dataAxi_rd_bits_last ? _GEN_733 : valid_3_5; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_863 = io_dataAxi_rd_bits_last ? _GEN_734 : valid_3_6; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_864 = io_dataAxi_rd_bits_last ? _GEN_735 : valid_3_7; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_865 = io_dataAxi_rd_bits_last ? _GEN_736 : valid_3_8; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_866 = io_dataAxi_rd_bits_last ? _GEN_737 : valid_3_9; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_867 = io_dataAxi_rd_bits_last ? _GEN_738 : valid_3_10; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_868 = io_dataAxi_rd_bits_last ? _GEN_739 : valid_3_11; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_869 = io_dataAxi_rd_bits_last ? _GEN_740 : valid_3_12; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_870 = io_dataAxi_rd_bits_last ? _GEN_741 : valid_3_13; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_871 = io_dataAxi_rd_bits_last ? _GEN_742 : valid_3_14; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire  _GEN_872 = io_dataAxi_rd_bits_last ? _GEN_743 : valid_3_15; // @[dcache.scala 272:46 dcache.scala 93:26]
  wire [2:0] _GEN_873 = io_dataAxi_rd_bits_last ? 3'h0 : state; // @[dcache.scala 272:46 dcache.scala 276:27 dcache.scala 153:24]
  wire [2:0] _GEN_874 = axiRdataEn & io_dataAxi_rd_valid ? _offset_T_1 : offset; // @[dcache.scala 265:52 dcache.scala 266:24 dcache.scala 111:34]
  wire [63:0] _GEN_876 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_615 : rdatabuf; // @[dcache.scala 265:52 dcache.scala 112:34]
  wire  _GEN_877 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_744 : axiRdataEn; // @[dcache.scala 265:52 dcache.scala 220:34]
  wire [21:0] _GEN_878 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_745 : tag_0_0; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_879 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_746 : tag_0_1; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_880 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_747 : tag_0_2; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_881 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_748 : tag_0_3; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_882 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_749 : tag_0_4; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_883 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_750 : tag_0_5; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_884 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_751 : tag_0_6; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_885 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_752 : tag_0_7; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_886 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_753 : tag_0_8; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_887 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_754 : tag_0_9; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_888 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_755 : tag_0_10; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_889 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_756 : tag_0_11; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_890 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_757 : tag_0_12; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_891 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_758 : tag_0_13; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_892 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_759 : tag_0_14; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_893 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_760 : tag_0_15; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_894 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_761 : tag_1_0; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_895 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_762 : tag_1_1; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_896 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_763 : tag_1_2; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_897 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_764 : tag_1_3; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_898 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_765 : tag_1_4; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_899 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_766 : tag_1_5; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_900 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_767 : tag_1_6; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_901 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_768 : tag_1_7; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_902 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_769 : tag_1_8; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_903 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_770 : tag_1_9; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_904 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_771 : tag_1_10; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_905 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_772 : tag_1_11; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_906 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_773 : tag_1_12; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_907 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_774 : tag_1_13; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_908 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_775 : tag_1_14; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_909 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_776 : tag_1_15; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_910 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_777 : tag_2_0; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_911 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_778 : tag_2_1; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_912 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_779 : tag_2_2; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_913 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_780 : tag_2_3; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_914 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_781 : tag_2_4; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_915 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_782 : tag_2_5; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_916 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_783 : tag_2_6; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_917 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_784 : tag_2_7; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_918 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_785 : tag_2_8; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_919 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_786 : tag_2_9; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_920 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_787 : tag_2_10; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_921 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_788 : tag_2_11; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_922 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_789 : tag_2_12; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_923 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_790 : tag_2_13; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_924 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_791 : tag_2_14; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_925 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_792 : tag_2_15; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_926 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_793 : tag_3_0; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_927 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_794 : tag_3_1; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_928 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_795 : tag_3_2; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_929 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_796 : tag_3_3; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_930 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_797 : tag_3_4; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_931 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_798 : tag_3_5; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_932 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_799 : tag_3_6; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_933 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_800 : tag_3_7; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_934 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_801 : tag_3_8; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_935 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_802 : tag_3_9; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_936 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_803 : tag_3_10; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_937 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_804 : tag_3_11; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_938 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_805 : tag_3_12; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_939 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_806 : tag_3_13; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_940 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_807 : tag_3_14; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire [21:0] _GEN_941 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_808 : tag_3_15; // @[dcache.scala 265:52 dcache.scala 92:26]
  wire  _GEN_942 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_809 : valid_0_0; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_943 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_810 : valid_0_1; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_944 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_811 : valid_0_2; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_945 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_812 : valid_0_3; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_946 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_813 : valid_0_4; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_947 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_814 : valid_0_5; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_948 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_815 : valid_0_6; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_949 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_816 : valid_0_7; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_950 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_817 : valid_0_8; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_951 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_818 : valid_0_9; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_952 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_819 : valid_0_10; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_953 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_820 : valid_0_11; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_954 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_821 : valid_0_12; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_955 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_822 : valid_0_13; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_956 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_823 : valid_0_14; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_957 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_824 : valid_0_15; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_958 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_825 : valid_1_0; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_959 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_826 : valid_1_1; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_960 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_827 : valid_1_2; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_961 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_828 : valid_1_3; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_962 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_829 : valid_1_4; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_963 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_830 : valid_1_5; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_964 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_831 : valid_1_6; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_965 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_832 : valid_1_7; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_966 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_833 : valid_1_8; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_967 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_834 : valid_1_9; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_968 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_835 : valid_1_10; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_969 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_836 : valid_1_11; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_970 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_837 : valid_1_12; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_971 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_838 : valid_1_13; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_972 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_839 : valid_1_14; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_973 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_840 : valid_1_15; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_974 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_841 : valid_2_0; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_975 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_842 : valid_2_1; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_976 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_843 : valid_2_2; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_977 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_844 : valid_2_3; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_978 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_845 : valid_2_4; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_979 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_846 : valid_2_5; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_980 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_847 : valid_2_6; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_981 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_848 : valid_2_7; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_982 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_849 : valid_2_8; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_983 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_850 : valid_2_9; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_984 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_851 : valid_2_10; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_985 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_852 : valid_2_11; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_986 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_853 : valid_2_12; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_987 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_854 : valid_2_13; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_988 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_855 : valid_2_14; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_989 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_856 : valid_2_15; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_990 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_857 : valid_3_0; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_991 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_858 : valid_3_1; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_992 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_859 : valid_3_2; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_993 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_860 : valid_3_3; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_994 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_861 : valid_3_4; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_995 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_862 : valid_3_5; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_996 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_863 : valid_3_6; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_997 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_864 : valid_3_7; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_998 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_865 : valid_3_8; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_999 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_866 : valid_3_9; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_1000 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_867 : valid_3_10; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_1001 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_868 : valid_3_11; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_1002 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_869 : valid_3_12; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_1003 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_870 : valid_3_13; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_1004 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_871 : valid_3_14; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire  _GEN_1005 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_872 : valid_3_15; // @[dcache.scala 265:52 dcache.scala 93:26]
  wire [2:0] _GEN_1006 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_873 : state; // @[dcache.scala 265:52 dcache.scala 153:24]
  wire [2:0] _GEN_1007 = axiWaddrEn & io_dataAxi_wa_ready ? 3'h4 : state; // @[dcache.scala 282:52 dcache.scala 283:29 dcache.scala 153:24]
  wire  _GEN_1008 = axiWaddrEn & io_dataAxi_wa_ready ? 1'h0 : axiWaddrEn; // @[dcache.scala 282:52 dcache.scala 284:29 dcache.scala 221:34]
  wire  _GEN_1009 = axiWaddrEn & io_dataAxi_wa_ready | axiWdataEn; // @[dcache.scala 282:52 dcache.scala 285:29 dcache.scala 224:34]
  wire  _GEN_1010 = _GEN_2695 & _GEN_2726 ? 1'h0 : valid_0_0; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1011 = _GEN_2695 & _GEN_2696 ? 1'h0 : valid_0_1; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1012 = _GEN_2695 & _GEN_2698 ? 1'h0 : valid_0_2; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1013 = _GEN_2695 & _GEN_2700 ? 1'h0 : valid_0_3; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1014 = _GEN_2695 & _GEN_2702 ? 1'h0 : valid_0_4; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1015 = _GEN_2695 & _GEN_2704 ? 1'h0 : valid_0_5; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1016 = _GEN_2695 & _GEN_2706 ? 1'h0 : valid_0_6; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1017 = _GEN_2695 & _GEN_2708 ? 1'h0 : valid_0_7; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1018 = _GEN_2695 & _GEN_2710 ? 1'h0 : valid_0_8; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1019 = _GEN_2695 & _GEN_2712 ? 1'h0 : valid_0_9; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1020 = _GEN_2695 & _GEN_2714 ? 1'h0 : valid_0_10; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1021 = _GEN_2695 & _GEN_2716 ? 1'h0 : valid_0_11; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1022 = _GEN_2695 & _GEN_2718 ? 1'h0 : valid_0_12; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1023 = _GEN_2695 & _GEN_2720 ? 1'h0 : valid_0_13; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1024 = _GEN_2695 & _GEN_2722 ? 1'h0 : valid_0_14; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1025 = _GEN_2695 & _GEN_2724 ? 1'h0 : valid_0_15; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1026 = _rdata128_T & _GEN_2726 ? 1'h0 : valid_1_0; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1027 = _rdata128_T & _GEN_2696 ? 1'h0 : valid_1_1; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1028 = _rdata128_T & _GEN_2698 ? 1'h0 : valid_1_2; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1029 = _rdata128_T & _GEN_2700 ? 1'h0 : valid_1_3; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1030 = _rdata128_T & _GEN_2702 ? 1'h0 : valid_1_4; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1031 = _rdata128_T & _GEN_2704 ? 1'h0 : valid_1_5; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1032 = _rdata128_T & _GEN_2706 ? 1'h0 : valid_1_6; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1033 = _rdata128_T & _GEN_2708 ? 1'h0 : valid_1_7; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1034 = _rdata128_T & _GEN_2710 ? 1'h0 : valid_1_8; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1035 = _rdata128_T & _GEN_2712 ? 1'h0 : valid_1_9; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1036 = _rdata128_T & _GEN_2714 ? 1'h0 : valid_1_10; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1037 = _rdata128_T & _GEN_2716 ? 1'h0 : valid_1_11; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1038 = _rdata128_T & _GEN_2718 ? 1'h0 : valid_1_12; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1039 = _rdata128_T & _GEN_2720 ? 1'h0 : valid_1_13; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1040 = _rdata128_T & _GEN_2722 ? 1'h0 : valid_1_14; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1041 = _rdata128_T & _GEN_2724 ? 1'h0 : valid_1_15; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1042 = _rdata128_T_2 & _GEN_2726 ? 1'h0 : valid_2_0; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1043 = _rdata128_T_2 & _GEN_2696 ? 1'h0 : valid_2_1; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1044 = _rdata128_T_2 & _GEN_2698 ? 1'h0 : valid_2_2; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1045 = _rdata128_T_2 & _GEN_2700 ? 1'h0 : valid_2_3; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1046 = _rdata128_T_2 & _GEN_2702 ? 1'h0 : valid_2_4; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1047 = _rdata128_T_2 & _GEN_2704 ? 1'h0 : valid_2_5; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1048 = _rdata128_T_2 & _GEN_2706 ? 1'h0 : valid_2_6; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1049 = _rdata128_T_2 & _GEN_2708 ? 1'h0 : valid_2_7; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1050 = _rdata128_T_2 & _GEN_2710 ? 1'h0 : valid_2_8; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1051 = _rdata128_T_2 & _GEN_2712 ? 1'h0 : valid_2_9; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1052 = _rdata128_T_2 & _GEN_2714 ? 1'h0 : valid_2_10; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1053 = _rdata128_T_2 & _GEN_2716 ? 1'h0 : valid_2_11; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1054 = _rdata128_T_2 & _GEN_2718 ? 1'h0 : valid_2_12; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1055 = _rdata128_T_2 & _GEN_2720 ? 1'h0 : valid_2_13; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1056 = _rdata128_T_2 & _GEN_2722 ? 1'h0 : valid_2_14; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1057 = _rdata128_T_2 & _GEN_2724 ? 1'h0 : valid_2_15; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1058 = _rdata128_T_4 & _GEN_2726 ? 1'h0 : valid_3_0; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1059 = _rdata128_T_4 & _GEN_2696 ? 1'h0 : valid_3_1; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1060 = _rdata128_T_4 & _GEN_2698 ? 1'h0 : valid_3_2; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1061 = _rdata128_T_4 & _GEN_2700 ? 1'h0 : valid_3_3; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1062 = _rdata128_T_4 & _GEN_2702 ? 1'h0 : valid_3_4; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1063 = _rdata128_T_4 & _GEN_2704 ? 1'h0 : valid_3_5; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1064 = _rdata128_T_4 & _GEN_2706 ? 1'h0 : valid_3_6; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1065 = _rdata128_T_4 & _GEN_2708 ? 1'h0 : valid_3_7; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1066 = _rdata128_T_4 & _GEN_2710 ? 1'h0 : valid_3_8; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1067 = _rdata128_T_4 & _GEN_2712 ? 1'h0 : valid_3_9; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1068 = _rdata128_T_4 & _GEN_2714 ? 1'h0 : valid_3_10; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1069 = _rdata128_T_4 & _GEN_2716 ? 1'h0 : valid_3_11; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1070 = _rdata128_T_4 & _GEN_2718 ? 1'h0 : valid_3_12; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1071 = _rdata128_T_4 & _GEN_2720 ? 1'h0 : valid_3_13; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1072 = _rdata128_T_4 & _GEN_2722 ? 1'h0 : valid_3_14; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1073 = _rdata128_T_4 & _GEN_2724 ? 1'h0 : valid_3_15; // @[dcache.scala 296:51 dcache.scala 296:51 dcache.scala 93:26]
  wire  _GEN_1074 = _GEN_2695 & _GEN_2726 ? 1'h0 : _GEN_390; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1075 = _GEN_2695 & _GEN_2696 ? 1'h0 : _GEN_391; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1076 = _GEN_2695 & _GEN_2698 ? 1'h0 : _GEN_392; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1077 = _GEN_2695 & _GEN_2700 ? 1'h0 : _GEN_393; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1078 = _GEN_2695 & _GEN_2702 ? 1'h0 : _GEN_394; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1079 = _GEN_2695 & _GEN_2704 ? 1'h0 : _GEN_395; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1080 = _GEN_2695 & _GEN_2706 ? 1'h0 : _GEN_396; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1081 = _GEN_2695 & _GEN_2708 ? 1'h0 : _GEN_397; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1082 = _GEN_2695 & _GEN_2710 ? 1'h0 : _GEN_398; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1083 = _GEN_2695 & _GEN_2712 ? 1'h0 : _GEN_399; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1084 = _GEN_2695 & _GEN_2714 ? 1'h0 : _GEN_400; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1085 = _GEN_2695 & _GEN_2716 ? 1'h0 : _GEN_401; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1086 = _GEN_2695 & _GEN_2718 ? 1'h0 : _GEN_402; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1087 = _GEN_2695 & _GEN_2720 ? 1'h0 : _GEN_403; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1088 = _GEN_2695 & _GEN_2722 ? 1'h0 : _GEN_404; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1089 = _GEN_2695 & _GEN_2724 ? 1'h0 : _GEN_405; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1090 = _rdata128_T & _GEN_2726 ? 1'h0 : _GEN_406; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1091 = _rdata128_T & _GEN_2696 ? 1'h0 : _GEN_407; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1092 = _rdata128_T & _GEN_2698 ? 1'h0 : _GEN_408; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1093 = _rdata128_T & _GEN_2700 ? 1'h0 : _GEN_409; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1094 = _rdata128_T & _GEN_2702 ? 1'h0 : _GEN_410; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1095 = _rdata128_T & _GEN_2704 ? 1'h0 : _GEN_411; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1096 = _rdata128_T & _GEN_2706 ? 1'h0 : _GEN_412; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1097 = _rdata128_T & _GEN_2708 ? 1'h0 : _GEN_413; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1098 = _rdata128_T & _GEN_2710 ? 1'h0 : _GEN_414; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1099 = _rdata128_T & _GEN_2712 ? 1'h0 : _GEN_415; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1100 = _rdata128_T & _GEN_2714 ? 1'h0 : _GEN_416; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1101 = _rdata128_T & _GEN_2716 ? 1'h0 : _GEN_417; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1102 = _rdata128_T & _GEN_2718 ? 1'h0 : _GEN_418; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1103 = _rdata128_T & _GEN_2720 ? 1'h0 : _GEN_419; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1104 = _rdata128_T & _GEN_2722 ? 1'h0 : _GEN_420; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1105 = _rdata128_T & _GEN_2724 ? 1'h0 : _GEN_421; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1106 = _rdata128_T_2 & _GEN_2726 ? 1'h0 : _GEN_422; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1107 = _rdata128_T_2 & _GEN_2696 ? 1'h0 : _GEN_423; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1108 = _rdata128_T_2 & _GEN_2698 ? 1'h0 : _GEN_424; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1109 = _rdata128_T_2 & _GEN_2700 ? 1'h0 : _GEN_425; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1110 = _rdata128_T_2 & _GEN_2702 ? 1'h0 : _GEN_426; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1111 = _rdata128_T_2 & _GEN_2704 ? 1'h0 : _GEN_427; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1112 = _rdata128_T_2 & _GEN_2706 ? 1'h0 : _GEN_428; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1113 = _rdata128_T_2 & _GEN_2708 ? 1'h0 : _GEN_429; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1114 = _rdata128_T_2 & _GEN_2710 ? 1'h0 : _GEN_430; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1115 = _rdata128_T_2 & _GEN_2712 ? 1'h0 : _GEN_431; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1116 = _rdata128_T_2 & _GEN_2714 ? 1'h0 : _GEN_432; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1117 = _rdata128_T_2 & _GEN_2716 ? 1'h0 : _GEN_433; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1118 = _rdata128_T_2 & _GEN_2718 ? 1'h0 : _GEN_434; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1119 = _rdata128_T_2 & _GEN_2720 ? 1'h0 : _GEN_435; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1120 = _rdata128_T_2 & _GEN_2722 ? 1'h0 : _GEN_436; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1121 = _rdata128_T_2 & _GEN_2724 ? 1'h0 : _GEN_437; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1122 = _rdata128_T_4 & _GEN_2726 ? 1'h0 : _GEN_438; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1123 = _rdata128_T_4 & _GEN_2696 ? 1'h0 : _GEN_439; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1124 = _rdata128_T_4 & _GEN_2698 ? 1'h0 : _GEN_440; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1125 = _rdata128_T_4 & _GEN_2700 ? 1'h0 : _GEN_441; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1126 = _rdata128_T_4 & _GEN_2702 ? 1'h0 : _GEN_442; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1127 = _rdata128_T_4 & _GEN_2704 ? 1'h0 : _GEN_443; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1128 = _rdata128_T_4 & _GEN_2706 ? 1'h0 : _GEN_444; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1129 = _rdata128_T_4 & _GEN_2708 ? 1'h0 : _GEN_445; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1130 = _rdata128_T_4 & _GEN_2710 ? 1'h0 : _GEN_446; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1131 = _rdata128_T_4 & _GEN_2712 ? 1'h0 : _GEN_447; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1132 = _rdata128_T_4 & _GEN_2714 ? 1'h0 : _GEN_448; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1133 = _rdata128_T_4 & _GEN_2716 ? 1'h0 : _GEN_449; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1134 = _rdata128_T_4 & _GEN_2718 ? 1'h0 : _GEN_450; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1135 = _rdata128_T_4 & _GEN_2720 ? 1'h0 : _GEN_451; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1136 = _rdata128_T_4 & _GEN_2722 ? 1'h0 : _GEN_452; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire  _GEN_1137 = _rdata128_T_4 & _GEN_2724 ? 1'h0 : _GEN_453; // @[dcache.scala 297:51 dcache.scala 297:51]
  wire [2:0] _GEN_1138 = io_dataAxi_wd_bits_last ? 3'h0 : state; // @[dcache.scala 293:46 dcache.scala 294:27 dcache.scala 153:24]
  wire  _GEN_1140 = io_dataAxi_wd_bits_last ? _GEN_1010 : valid_0_0; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1141 = io_dataAxi_wd_bits_last ? _GEN_1011 : valid_0_1; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1142 = io_dataAxi_wd_bits_last ? _GEN_1012 : valid_0_2; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1143 = io_dataAxi_wd_bits_last ? _GEN_1013 : valid_0_3; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1144 = io_dataAxi_wd_bits_last ? _GEN_1014 : valid_0_4; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1145 = io_dataAxi_wd_bits_last ? _GEN_1015 : valid_0_5; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1146 = io_dataAxi_wd_bits_last ? _GEN_1016 : valid_0_6; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1147 = io_dataAxi_wd_bits_last ? _GEN_1017 : valid_0_7; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1148 = io_dataAxi_wd_bits_last ? _GEN_1018 : valid_0_8; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1149 = io_dataAxi_wd_bits_last ? _GEN_1019 : valid_0_9; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1150 = io_dataAxi_wd_bits_last ? _GEN_1020 : valid_0_10; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1151 = io_dataAxi_wd_bits_last ? _GEN_1021 : valid_0_11; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1152 = io_dataAxi_wd_bits_last ? _GEN_1022 : valid_0_12; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1153 = io_dataAxi_wd_bits_last ? _GEN_1023 : valid_0_13; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1154 = io_dataAxi_wd_bits_last ? _GEN_1024 : valid_0_14; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1155 = io_dataAxi_wd_bits_last ? _GEN_1025 : valid_0_15; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1156 = io_dataAxi_wd_bits_last ? _GEN_1026 : valid_1_0; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1157 = io_dataAxi_wd_bits_last ? _GEN_1027 : valid_1_1; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1158 = io_dataAxi_wd_bits_last ? _GEN_1028 : valid_1_2; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1159 = io_dataAxi_wd_bits_last ? _GEN_1029 : valid_1_3; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1160 = io_dataAxi_wd_bits_last ? _GEN_1030 : valid_1_4; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1161 = io_dataAxi_wd_bits_last ? _GEN_1031 : valid_1_5; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1162 = io_dataAxi_wd_bits_last ? _GEN_1032 : valid_1_6; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1163 = io_dataAxi_wd_bits_last ? _GEN_1033 : valid_1_7; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1164 = io_dataAxi_wd_bits_last ? _GEN_1034 : valid_1_8; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1165 = io_dataAxi_wd_bits_last ? _GEN_1035 : valid_1_9; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1166 = io_dataAxi_wd_bits_last ? _GEN_1036 : valid_1_10; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1167 = io_dataAxi_wd_bits_last ? _GEN_1037 : valid_1_11; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1168 = io_dataAxi_wd_bits_last ? _GEN_1038 : valid_1_12; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1169 = io_dataAxi_wd_bits_last ? _GEN_1039 : valid_1_13; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1170 = io_dataAxi_wd_bits_last ? _GEN_1040 : valid_1_14; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1171 = io_dataAxi_wd_bits_last ? _GEN_1041 : valid_1_15; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1172 = io_dataAxi_wd_bits_last ? _GEN_1042 : valid_2_0; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1173 = io_dataAxi_wd_bits_last ? _GEN_1043 : valid_2_1; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1174 = io_dataAxi_wd_bits_last ? _GEN_1044 : valid_2_2; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1175 = io_dataAxi_wd_bits_last ? _GEN_1045 : valid_2_3; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1176 = io_dataAxi_wd_bits_last ? _GEN_1046 : valid_2_4; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1177 = io_dataAxi_wd_bits_last ? _GEN_1047 : valid_2_5; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1178 = io_dataAxi_wd_bits_last ? _GEN_1048 : valid_2_6; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1179 = io_dataAxi_wd_bits_last ? _GEN_1049 : valid_2_7; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1180 = io_dataAxi_wd_bits_last ? _GEN_1050 : valid_2_8; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1181 = io_dataAxi_wd_bits_last ? _GEN_1051 : valid_2_9; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1182 = io_dataAxi_wd_bits_last ? _GEN_1052 : valid_2_10; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1183 = io_dataAxi_wd_bits_last ? _GEN_1053 : valid_2_11; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1184 = io_dataAxi_wd_bits_last ? _GEN_1054 : valid_2_12; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1185 = io_dataAxi_wd_bits_last ? _GEN_1055 : valid_2_13; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1186 = io_dataAxi_wd_bits_last ? _GEN_1056 : valid_2_14; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1187 = io_dataAxi_wd_bits_last ? _GEN_1057 : valid_2_15; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1188 = io_dataAxi_wd_bits_last ? _GEN_1058 : valid_3_0; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1189 = io_dataAxi_wd_bits_last ? _GEN_1059 : valid_3_1; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1190 = io_dataAxi_wd_bits_last ? _GEN_1060 : valid_3_2; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1191 = io_dataAxi_wd_bits_last ? _GEN_1061 : valid_3_3; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1192 = io_dataAxi_wd_bits_last ? _GEN_1062 : valid_3_4; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1193 = io_dataAxi_wd_bits_last ? _GEN_1063 : valid_3_5; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1194 = io_dataAxi_wd_bits_last ? _GEN_1064 : valid_3_6; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1195 = io_dataAxi_wd_bits_last ? _GEN_1065 : valid_3_7; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1196 = io_dataAxi_wd_bits_last ? _GEN_1066 : valid_3_8; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1197 = io_dataAxi_wd_bits_last ? _GEN_1067 : valid_3_9; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1198 = io_dataAxi_wd_bits_last ? _GEN_1068 : valid_3_10; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1199 = io_dataAxi_wd_bits_last ? _GEN_1069 : valid_3_11; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1200 = io_dataAxi_wd_bits_last ? _GEN_1070 : valid_3_12; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1201 = io_dataAxi_wd_bits_last ? _GEN_1071 : valid_3_13; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1202 = io_dataAxi_wd_bits_last ? _GEN_1072 : valid_3_14; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1203 = io_dataAxi_wd_bits_last ? _GEN_1073 : valid_3_15; // @[dcache.scala 293:46 dcache.scala 93:26]
  wire  _GEN_1204 = io_dataAxi_wd_bits_last ? _GEN_1074 : _GEN_390; // @[dcache.scala 293:46]
  wire  _GEN_1205 = io_dataAxi_wd_bits_last ? _GEN_1075 : _GEN_391; // @[dcache.scala 293:46]
  wire  _GEN_1206 = io_dataAxi_wd_bits_last ? _GEN_1076 : _GEN_392; // @[dcache.scala 293:46]
  wire  _GEN_1207 = io_dataAxi_wd_bits_last ? _GEN_1077 : _GEN_393; // @[dcache.scala 293:46]
  wire  _GEN_1208 = io_dataAxi_wd_bits_last ? _GEN_1078 : _GEN_394; // @[dcache.scala 293:46]
  wire  _GEN_1209 = io_dataAxi_wd_bits_last ? _GEN_1079 : _GEN_395; // @[dcache.scala 293:46]
  wire  _GEN_1210 = io_dataAxi_wd_bits_last ? _GEN_1080 : _GEN_396; // @[dcache.scala 293:46]
  wire  _GEN_1211 = io_dataAxi_wd_bits_last ? _GEN_1081 : _GEN_397; // @[dcache.scala 293:46]
  wire  _GEN_1212 = io_dataAxi_wd_bits_last ? _GEN_1082 : _GEN_398; // @[dcache.scala 293:46]
  wire  _GEN_1213 = io_dataAxi_wd_bits_last ? _GEN_1083 : _GEN_399; // @[dcache.scala 293:46]
  wire  _GEN_1214 = io_dataAxi_wd_bits_last ? _GEN_1084 : _GEN_400; // @[dcache.scala 293:46]
  wire  _GEN_1215 = io_dataAxi_wd_bits_last ? _GEN_1085 : _GEN_401; // @[dcache.scala 293:46]
  wire  _GEN_1216 = io_dataAxi_wd_bits_last ? _GEN_1086 : _GEN_402; // @[dcache.scala 293:46]
  wire  _GEN_1217 = io_dataAxi_wd_bits_last ? _GEN_1087 : _GEN_403; // @[dcache.scala 293:46]
  wire  _GEN_1218 = io_dataAxi_wd_bits_last ? _GEN_1088 : _GEN_404; // @[dcache.scala 293:46]
  wire  _GEN_1219 = io_dataAxi_wd_bits_last ? _GEN_1089 : _GEN_405; // @[dcache.scala 293:46]
  wire  _GEN_1220 = io_dataAxi_wd_bits_last ? _GEN_1090 : _GEN_406; // @[dcache.scala 293:46]
  wire  _GEN_1221 = io_dataAxi_wd_bits_last ? _GEN_1091 : _GEN_407; // @[dcache.scala 293:46]
  wire  _GEN_1222 = io_dataAxi_wd_bits_last ? _GEN_1092 : _GEN_408; // @[dcache.scala 293:46]
  wire  _GEN_1223 = io_dataAxi_wd_bits_last ? _GEN_1093 : _GEN_409; // @[dcache.scala 293:46]
  wire  _GEN_1224 = io_dataAxi_wd_bits_last ? _GEN_1094 : _GEN_410; // @[dcache.scala 293:46]
  wire  _GEN_1225 = io_dataAxi_wd_bits_last ? _GEN_1095 : _GEN_411; // @[dcache.scala 293:46]
  wire  _GEN_1226 = io_dataAxi_wd_bits_last ? _GEN_1096 : _GEN_412; // @[dcache.scala 293:46]
  wire  _GEN_1227 = io_dataAxi_wd_bits_last ? _GEN_1097 : _GEN_413; // @[dcache.scala 293:46]
  wire  _GEN_1228 = io_dataAxi_wd_bits_last ? _GEN_1098 : _GEN_414; // @[dcache.scala 293:46]
  wire  _GEN_1229 = io_dataAxi_wd_bits_last ? _GEN_1099 : _GEN_415; // @[dcache.scala 293:46]
  wire  _GEN_1230 = io_dataAxi_wd_bits_last ? _GEN_1100 : _GEN_416; // @[dcache.scala 293:46]
  wire  _GEN_1231 = io_dataAxi_wd_bits_last ? _GEN_1101 : _GEN_417; // @[dcache.scala 293:46]
  wire  _GEN_1232 = io_dataAxi_wd_bits_last ? _GEN_1102 : _GEN_418; // @[dcache.scala 293:46]
  wire  _GEN_1233 = io_dataAxi_wd_bits_last ? _GEN_1103 : _GEN_419; // @[dcache.scala 293:46]
  wire  _GEN_1234 = io_dataAxi_wd_bits_last ? _GEN_1104 : _GEN_420; // @[dcache.scala 293:46]
  wire  _GEN_1235 = io_dataAxi_wd_bits_last ? _GEN_1105 : _GEN_421; // @[dcache.scala 293:46]
  wire  _GEN_1236 = io_dataAxi_wd_bits_last ? _GEN_1106 : _GEN_422; // @[dcache.scala 293:46]
  wire  _GEN_1237 = io_dataAxi_wd_bits_last ? _GEN_1107 : _GEN_423; // @[dcache.scala 293:46]
  wire  _GEN_1238 = io_dataAxi_wd_bits_last ? _GEN_1108 : _GEN_424; // @[dcache.scala 293:46]
  wire  _GEN_1239 = io_dataAxi_wd_bits_last ? _GEN_1109 : _GEN_425; // @[dcache.scala 293:46]
  wire  _GEN_1240 = io_dataAxi_wd_bits_last ? _GEN_1110 : _GEN_426; // @[dcache.scala 293:46]
  wire  _GEN_1241 = io_dataAxi_wd_bits_last ? _GEN_1111 : _GEN_427; // @[dcache.scala 293:46]
  wire  _GEN_1242 = io_dataAxi_wd_bits_last ? _GEN_1112 : _GEN_428; // @[dcache.scala 293:46]
  wire  _GEN_1243 = io_dataAxi_wd_bits_last ? _GEN_1113 : _GEN_429; // @[dcache.scala 293:46]
  wire  _GEN_1244 = io_dataAxi_wd_bits_last ? _GEN_1114 : _GEN_430; // @[dcache.scala 293:46]
  wire  _GEN_1245 = io_dataAxi_wd_bits_last ? _GEN_1115 : _GEN_431; // @[dcache.scala 293:46]
  wire  _GEN_1246 = io_dataAxi_wd_bits_last ? _GEN_1116 : _GEN_432; // @[dcache.scala 293:46]
  wire  _GEN_1247 = io_dataAxi_wd_bits_last ? _GEN_1117 : _GEN_433; // @[dcache.scala 293:46]
  wire  _GEN_1248 = io_dataAxi_wd_bits_last ? _GEN_1118 : _GEN_434; // @[dcache.scala 293:46]
  wire  _GEN_1249 = io_dataAxi_wd_bits_last ? _GEN_1119 : _GEN_435; // @[dcache.scala 293:46]
  wire  _GEN_1250 = io_dataAxi_wd_bits_last ? _GEN_1120 : _GEN_436; // @[dcache.scala 293:46]
  wire  _GEN_1251 = io_dataAxi_wd_bits_last ? _GEN_1121 : _GEN_437; // @[dcache.scala 293:46]
  wire  _GEN_1252 = io_dataAxi_wd_bits_last ? _GEN_1122 : _GEN_438; // @[dcache.scala 293:46]
  wire  _GEN_1253 = io_dataAxi_wd_bits_last ? _GEN_1123 : _GEN_439; // @[dcache.scala 293:46]
  wire  _GEN_1254 = io_dataAxi_wd_bits_last ? _GEN_1124 : _GEN_440; // @[dcache.scala 293:46]
  wire  _GEN_1255 = io_dataAxi_wd_bits_last ? _GEN_1125 : _GEN_441; // @[dcache.scala 293:46]
  wire  _GEN_1256 = io_dataAxi_wd_bits_last ? _GEN_1126 : _GEN_442; // @[dcache.scala 293:46]
  wire  _GEN_1257 = io_dataAxi_wd_bits_last ? _GEN_1127 : _GEN_443; // @[dcache.scala 293:46]
  wire  _GEN_1258 = io_dataAxi_wd_bits_last ? _GEN_1128 : _GEN_444; // @[dcache.scala 293:46]
  wire  _GEN_1259 = io_dataAxi_wd_bits_last ? _GEN_1129 : _GEN_445; // @[dcache.scala 293:46]
  wire  _GEN_1260 = io_dataAxi_wd_bits_last ? _GEN_1130 : _GEN_446; // @[dcache.scala 293:46]
  wire  _GEN_1261 = io_dataAxi_wd_bits_last ? _GEN_1131 : _GEN_447; // @[dcache.scala 293:46]
  wire  _GEN_1262 = io_dataAxi_wd_bits_last ? _GEN_1132 : _GEN_448; // @[dcache.scala 293:46]
  wire  _GEN_1263 = io_dataAxi_wd_bits_last ? _GEN_1133 : _GEN_449; // @[dcache.scala 293:46]
  wire  _GEN_1264 = io_dataAxi_wd_bits_last ? _GEN_1134 : _GEN_450; // @[dcache.scala 293:46]
  wire  _GEN_1265 = io_dataAxi_wd_bits_last ? _GEN_1135 : _GEN_451; // @[dcache.scala 293:46]
  wire  _GEN_1266 = io_dataAxi_wd_bits_last ? _GEN_1136 : _GEN_452; // @[dcache.scala 293:46]
  wire  _GEN_1267 = io_dataAxi_wd_bits_last ? _GEN_1137 : _GEN_453; // @[dcache.scala 293:46]
  wire [2:0] _GEN_1268 = axiWdataEn & io_dataAxi_wd_ready ? _offset_T_1 : offset; // @[dcache.scala 290:52 dcache.scala 291:24 dcache.scala 111:34]
  wire  _GEN_1269 = axiWdataEn & io_dataAxi_wd_ready ? 1'h0 : 1'h1; // @[dcache.scala 290:52 dcache.scala 289:24]
  wire [2:0] _GEN_1270 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1138 : state; // @[dcache.scala 290:52 dcache.scala 153:24]
  wire  _GEN_1271 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1140 : valid_0_0; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1272 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1141 : valid_0_1; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1273 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1142 : valid_0_2; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1274 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1143 : valid_0_3; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1275 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1144 : valid_0_4; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1276 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1145 : valid_0_5; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1277 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1146 : valid_0_6; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1278 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1147 : valid_0_7; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1279 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1148 : valid_0_8; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1280 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1149 : valid_0_9; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1281 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1150 : valid_0_10; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1282 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1151 : valid_0_11; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1283 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1152 : valid_0_12; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1284 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1153 : valid_0_13; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1285 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1154 : valid_0_14; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1286 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1155 : valid_0_15; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1287 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1156 : valid_1_0; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1288 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1157 : valid_1_1; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1289 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1158 : valid_1_2; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1290 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1159 : valid_1_3; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1291 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1160 : valid_1_4; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1292 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1161 : valid_1_5; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1293 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1162 : valid_1_6; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1294 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1163 : valid_1_7; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1295 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1164 : valid_1_8; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1296 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1165 : valid_1_9; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1297 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1166 : valid_1_10; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1298 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1167 : valid_1_11; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1299 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1168 : valid_1_12; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1300 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1169 : valid_1_13; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1301 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1170 : valid_1_14; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1302 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1171 : valid_1_15; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1303 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1172 : valid_2_0; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1304 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1173 : valid_2_1; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1305 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1174 : valid_2_2; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1306 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1175 : valid_2_3; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1307 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1176 : valid_2_4; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1308 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1177 : valid_2_5; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1309 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1178 : valid_2_6; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1310 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1179 : valid_2_7; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1311 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1180 : valid_2_8; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1312 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1181 : valid_2_9; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1313 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1182 : valid_2_10; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1314 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1183 : valid_2_11; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1315 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1184 : valid_2_12; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1316 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1185 : valid_2_13; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1317 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1186 : valid_2_14; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1318 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1187 : valid_2_15; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1319 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1188 : valid_3_0; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1320 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1189 : valid_3_1; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1321 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1190 : valid_3_2; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1322 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1191 : valid_3_3; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1323 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1192 : valid_3_4; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1324 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1193 : valid_3_5; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1325 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1194 : valid_3_6; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1326 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1195 : valid_3_7; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1327 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1196 : valid_3_8; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1328 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1197 : valid_3_9; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1329 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1198 : valid_3_10; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1330 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1199 : valid_3_11; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1331 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1200 : valid_3_12; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1332 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1201 : valid_3_13; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1333 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1202 : valid_3_14; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1334 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1203 : valid_3_15; // @[dcache.scala 290:52 dcache.scala 93:26]
  wire  _GEN_1335 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1204 : _GEN_390; // @[dcache.scala 290:52]
  wire  _GEN_1336 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1205 : _GEN_391; // @[dcache.scala 290:52]
  wire  _GEN_1337 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1206 : _GEN_392; // @[dcache.scala 290:52]
  wire  _GEN_1338 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1207 : _GEN_393; // @[dcache.scala 290:52]
  wire  _GEN_1339 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1208 : _GEN_394; // @[dcache.scala 290:52]
  wire  _GEN_1340 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1209 : _GEN_395; // @[dcache.scala 290:52]
  wire  _GEN_1341 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1210 : _GEN_396; // @[dcache.scala 290:52]
  wire  _GEN_1342 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1211 : _GEN_397; // @[dcache.scala 290:52]
  wire  _GEN_1343 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1212 : _GEN_398; // @[dcache.scala 290:52]
  wire  _GEN_1344 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1213 : _GEN_399; // @[dcache.scala 290:52]
  wire  _GEN_1345 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1214 : _GEN_400; // @[dcache.scala 290:52]
  wire  _GEN_1346 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1215 : _GEN_401; // @[dcache.scala 290:52]
  wire  _GEN_1347 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1216 : _GEN_402; // @[dcache.scala 290:52]
  wire  _GEN_1348 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1217 : _GEN_403; // @[dcache.scala 290:52]
  wire  _GEN_1349 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1218 : _GEN_404; // @[dcache.scala 290:52]
  wire  _GEN_1350 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1219 : _GEN_405; // @[dcache.scala 290:52]
  wire  _GEN_1351 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1220 : _GEN_406; // @[dcache.scala 290:52]
  wire  _GEN_1352 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1221 : _GEN_407; // @[dcache.scala 290:52]
  wire  _GEN_1353 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1222 : _GEN_408; // @[dcache.scala 290:52]
  wire  _GEN_1354 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1223 : _GEN_409; // @[dcache.scala 290:52]
  wire  _GEN_1355 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1224 : _GEN_410; // @[dcache.scala 290:52]
  wire  _GEN_1356 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1225 : _GEN_411; // @[dcache.scala 290:52]
  wire  _GEN_1357 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1226 : _GEN_412; // @[dcache.scala 290:52]
  wire  _GEN_1358 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1227 : _GEN_413; // @[dcache.scala 290:52]
  wire  _GEN_1359 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1228 : _GEN_414; // @[dcache.scala 290:52]
  wire  _GEN_1360 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1229 : _GEN_415; // @[dcache.scala 290:52]
  wire  _GEN_1361 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1230 : _GEN_416; // @[dcache.scala 290:52]
  wire  _GEN_1362 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1231 : _GEN_417; // @[dcache.scala 290:52]
  wire  _GEN_1363 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1232 : _GEN_418; // @[dcache.scala 290:52]
  wire  _GEN_1364 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1233 : _GEN_419; // @[dcache.scala 290:52]
  wire  _GEN_1365 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1234 : _GEN_420; // @[dcache.scala 290:52]
  wire  _GEN_1366 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1235 : _GEN_421; // @[dcache.scala 290:52]
  wire  _GEN_1367 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1236 : _GEN_422; // @[dcache.scala 290:52]
  wire  _GEN_1368 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1237 : _GEN_423; // @[dcache.scala 290:52]
  wire  _GEN_1369 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1238 : _GEN_424; // @[dcache.scala 290:52]
  wire  _GEN_1370 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1239 : _GEN_425; // @[dcache.scala 290:52]
  wire  _GEN_1371 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1240 : _GEN_426; // @[dcache.scala 290:52]
  wire  _GEN_1372 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1241 : _GEN_427; // @[dcache.scala 290:52]
  wire  _GEN_1373 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1242 : _GEN_428; // @[dcache.scala 290:52]
  wire  _GEN_1374 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1243 : _GEN_429; // @[dcache.scala 290:52]
  wire  _GEN_1375 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1244 : _GEN_430; // @[dcache.scala 290:52]
  wire  _GEN_1376 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1245 : _GEN_431; // @[dcache.scala 290:52]
  wire  _GEN_1377 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1246 : _GEN_432; // @[dcache.scala 290:52]
  wire  _GEN_1378 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1247 : _GEN_433; // @[dcache.scala 290:52]
  wire  _GEN_1379 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1248 : _GEN_434; // @[dcache.scala 290:52]
  wire  _GEN_1380 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1249 : _GEN_435; // @[dcache.scala 290:52]
  wire  _GEN_1381 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1250 : _GEN_436; // @[dcache.scala 290:52]
  wire  _GEN_1382 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1251 : _GEN_437; // @[dcache.scala 290:52]
  wire  _GEN_1383 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1252 : _GEN_438; // @[dcache.scala 290:52]
  wire  _GEN_1384 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1253 : _GEN_439; // @[dcache.scala 290:52]
  wire  _GEN_1385 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1254 : _GEN_440; // @[dcache.scala 290:52]
  wire  _GEN_1386 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1255 : _GEN_441; // @[dcache.scala 290:52]
  wire  _GEN_1387 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1256 : _GEN_442; // @[dcache.scala 290:52]
  wire  _GEN_1388 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1257 : _GEN_443; // @[dcache.scala 290:52]
  wire  _GEN_1389 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1258 : _GEN_444; // @[dcache.scala 290:52]
  wire  _GEN_1390 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1259 : _GEN_445; // @[dcache.scala 290:52]
  wire  _GEN_1391 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1260 : _GEN_446; // @[dcache.scala 290:52]
  wire  _GEN_1392 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1261 : _GEN_447; // @[dcache.scala 290:52]
  wire  _GEN_1393 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1262 : _GEN_448; // @[dcache.scala 290:52]
  wire  _GEN_1394 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1263 : _GEN_449; // @[dcache.scala 290:52]
  wire  _GEN_1395 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1264 : _GEN_450; // @[dcache.scala 290:52]
  wire  _GEN_1396 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1265 : _GEN_451; // @[dcache.scala 290:52]
  wire  _GEN_1397 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1266 : _GEN_452; // @[dcache.scala 290:52]
  wire  _GEN_1398 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1267 : _GEN_453; // @[dcache.scala 290:52]
  wire  _T_84 = 3'h6 == state; // @[Conditional.scala 37:30]
  wire  _GEN_1399 = flush_done ? 1'h0 : _GEN_134; // @[dcache.scala 308:29 dcache.scala 309:25]
  wire [2:0] _GEN_1400 = flush_done ? 3'h0 : 3'h3; // @[dcache.scala 308:29 dcache.scala 310:23 dcache.scala 313:23]
  wire  _GEN_1401 = flush_done ? 1'h0 : valid_0_0; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1402 = flush_done ? 1'h0 : valid_0_1; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1403 = flush_done ? 1'h0 : valid_0_2; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1404 = flush_done ? 1'h0 : valid_0_3; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1405 = flush_done ? 1'h0 : valid_0_4; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1406 = flush_done ? 1'h0 : valid_0_5; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1407 = flush_done ? 1'h0 : valid_0_6; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1408 = flush_done ? 1'h0 : valid_0_7; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1409 = flush_done ? 1'h0 : valid_0_8; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1410 = flush_done ? 1'h0 : valid_0_9; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1411 = flush_done ? 1'h0 : valid_0_10; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1412 = flush_done ? 1'h0 : valid_0_11; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1413 = flush_done ? 1'h0 : valid_0_12; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1414 = flush_done ? 1'h0 : valid_0_13; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1415 = flush_done ? 1'h0 : valid_0_14; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1416 = flush_done ? 1'h0 : valid_0_15; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1417 = flush_done ? 1'h0 : valid_1_0; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1418 = flush_done ? 1'h0 : valid_1_1; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1419 = flush_done ? 1'h0 : valid_1_2; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1420 = flush_done ? 1'h0 : valid_1_3; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1421 = flush_done ? 1'h0 : valid_1_4; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1422 = flush_done ? 1'h0 : valid_1_5; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1423 = flush_done ? 1'h0 : valid_1_6; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1424 = flush_done ? 1'h0 : valid_1_7; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1425 = flush_done ? 1'h0 : valid_1_8; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1426 = flush_done ? 1'h0 : valid_1_9; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1427 = flush_done ? 1'h0 : valid_1_10; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1428 = flush_done ? 1'h0 : valid_1_11; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1429 = flush_done ? 1'h0 : valid_1_12; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1430 = flush_done ? 1'h0 : valid_1_13; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1431 = flush_done ? 1'h0 : valid_1_14; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1432 = flush_done ? 1'h0 : valid_1_15; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1433 = flush_done ? 1'h0 : valid_2_0; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1434 = flush_done ? 1'h0 : valid_2_1; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1435 = flush_done ? 1'h0 : valid_2_2; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1436 = flush_done ? 1'h0 : valid_2_3; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1437 = flush_done ? 1'h0 : valid_2_4; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1438 = flush_done ? 1'h0 : valid_2_5; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1439 = flush_done ? 1'h0 : valid_2_6; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1440 = flush_done ? 1'h0 : valid_2_7; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1441 = flush_done ? 1'h0 : valid_2_8; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1442 = flush_done ? 1'h0 : valid_2_9; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1443 = flush_done ? 1'h0 : valid_2_10; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1444 = flush_done ? 1'h0 : valid_2_11; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1445 = flush_done ? 1'h0 : valid_2_12; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1446 = flush_done ? 1'h0 : valid_2_13; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1447 = flush_done ? 1'h0 : valid_2_14; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1448 = flush_done ? 1'h0 : valid_2_15; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1449 = flush_done ? 1'h0 : valid_3_0; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1450 = flush_done ? 1'h0 : valid_3_1; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1451 = flush_done ? 1'h0 : valid_3_2; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1452 = flush_done ? 1'h0 : valid_3_3; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1453 = flush_done ? 1'h0 : valid_3_4; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1454 = flush_done ? 1'h0 : valid_3_5; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1455 = flush_done ? 1'h0 : valid_3_6; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1456 = flush_done ? 1'h0 : valid_3_7; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1457 = flush_done ? 1'h0 : valid_3_8; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1458 = flush_done ? 1'h0 : valid_3_9; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1459 = flush_done ? 1'h0 : valid_3_10; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1460 = flush_done ? 1'h0 : valid_3_11; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1461 = flush_done ? 1'h0 : valid_3_12; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1462 = flush_done ? 1'h0 : valid_3_13; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1463 = flush_done ? 1'h0 : valid_3_14; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1464 = flush_done ? 1'h0 : valid_3_15; // @[dcache.scala 308:29 dcache.scala 311:23 dcache.scala 93:26]
  wire  _GEN_1465 = flush_done ? axiWaddrEn : 1'h1; // @[dcache.scala 308:29 dcache.scala 221:34 dcache.scala 314:28]
  wire [1:0] _GEN_1466 = flush_done ? _GEN_129 : flush_way; // @[dcache.scala 308:29 dcache.scala 315:28]
  wire [3:0] _GEN_1467 = flush_done ? _GEN_133 : flush_idx; // @[dcache.scala 308:29 dcache.scala 316:28]
  wire  _GEN_1468 = _T_84 ? _GEN_1399 : _GEN_134; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_1469 = _T_84 ? _GEN_1400 : state; // @[Conditional.scala 39:67 dcache.scala 153:24]
  wire  _GEN_1470 = _T_84 ? _GEN_1401 : valid_0_0; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1471 = _T_84 ? _GEN_1402 : valid_0_1; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1472 = _T_84 ? _GEN_1403 : valid_0_2; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1473 = _T_84 ? _GEN_1404 : valid_0_3; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1474 = _T_84 ? _GEN_1405 : valid_0_4; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1475 = _T_84 ? _GEN_1406 : valid_0_5; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1476 = _T_84 ? _GEN_1407 : valid_0_6; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1477 = _T_84 ? _GEN_1408 : valid_0_7; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1478 = _T_84 ? _GEN_1409 : valid_0_8; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1479 = _T_84 ? _GEN_1410 : valid_0_9; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1480 = _T_84 ? _GEN_1411 : valid_0_10; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1481 = _T_84 ? _GEN_1412 : valid_0_11; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1482 = _T_84 ? _GEN_1413 : valid_0_12; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1483 = _T_84 ? _GEN_1414 : valid_0_13; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1484 = _T_84 ? _GEN_1415 : valid_0_14; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1485 = _T_84 ? _GEN_1416 : valid_0_15; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1486 = _T_84 ? _GEN_1417 : valid_1_0; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1487 = _T_84 ? _GEN_1418 : valid_1_1; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1488 = _T_84 ? _GEN_1419 : valid_1_2; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1489 = _T_84 ? _GEN_1420 : valid_1_3; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1490 = _T_84 ? _GEN_1421 : valid_1_4; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1491 = _T_84 ? _GEN_1422 : valid_1_5; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1492 = _T_84 ? _GEN_1423 : valid_1_6; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1493 = _T_84 ? _GEN_1424 : valid_1_7; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1494 = _T_84 ? _GEN_1425 : valid_1_8; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1495 = _T_84 ? _GEN_1426 : valid_1_9; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1496 = _T_84 ? _GEN_1427 : valid_1_10; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1497 = _T_84 ? _GEN_1428 : valid_1_11; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1498 = _T_84 ? _GEN_1429 : valid_1_12; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1499 = _T_84 ? _GEN_1430 : valid_1_13; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1500 = _T_84 ? _GEN_1431 : valid_1_14; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1501 = _T_84 ? _GEN_1432 : valid_1_15; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1502 = _T_84 ? _GEN_1433 : valid_2_0; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1503 = _T_84 ? _GEN_1434 : valid_2_1; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1504 = _T_84 ? _GEN_1435 : valid_2_2; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1505 = _T_84 ? _GEN_1436 : valid_2_3; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1506 = _T_84 ? _GEN_1437 : valid_2_4; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1507 = _T_84 ? _GEN_1438 : valid_2_5; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1508 = _T_84 ? _GEN_1439 : valid_2_6; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1509 = _T_84 ? _GEN_1440 : valid_2_7; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1510 = _T_84 ? _GEN_1441 : valid_2_8; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1511 = _T_84 ? _GEN_1442 : valid_2_9; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1512 = _T_84 ? _GEN_1443 : valid_2_10; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1513 = _T_84 ? _GEN_1444 : valid_2_11; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1514 = _T_84 ? _GEN_1445 : valid_2_12; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1515 = _T_84 ? _GEN_1446 : valid_2_13; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1516 = _T_84 ? _GEN_1447 : valid_2_14; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1517 = _T_84 ? _GEN_1448 : valid_2_15; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1518 = _T_84 ? _GEN_1449 : valid_3_0; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1519 = _T_84 ? _GEN_1450 : valid_3_1; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1520 = _T_84 ? _GEN_1451 : valid_3_2; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1521 = _T_84 ? _GEN_1452 : valid_3_3; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1522 = _T_84 ? _GEN_1453 : valid_3_4; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1523 = _T_84 ? _GEN_1454 : valid_3_5; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1524 = _T_84 ? _GEN_1455 : valid_3_6; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1525 = _T_84 ? _GEN_1456 : valid_3_7; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1526 = _T_84 ? _GEN_1457 : valid_3_8; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1527 = _T_84 ? _GEN_1458 : valid_3_9; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1528 = _T_84 ? _GEN_1459 : valid_3_10; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1529 = _T_84 ? _GEN_1460 : valid_3_11; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1530 = _T_84 ? _GEN_1461 : valid_3_12; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1531 = _T_84 ? _GEN_1462 : valid_3_13; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1532 = _T_84 ? _GEN_1463 : valid_3_14; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1533 = _T_84 ? _GEN_1464 : valid_3_15; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1534 = _T_84 ? _GEN_1465 : axiWaddrEn; // @[Conditional.scala 39:67 dcache.scala 221:34]
  wire [1:0] _GEN_1535 = _T_84 ? _GEN_1466 : _GEN_129; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_1536 = _T_84 ? _GEN_1467 : _GEN_133; // @[Conditional.scala 39:67]
  wire  _GEN_1539 = _T_83 ? 1'h0 : wait_r; // @[Conditional.scala 39:67 dcache.scala 304:21 dcache.scala 96:30]
  wire [2:0] _GEN_1540 = _T_83 ? 3'h0 : _GEN_1469; // @[Conditional.scala 39:67 dcache.scala 305:21]
  wire  _GEN_1541 = _T_83 ? _GEN_134 : _GEN_1468; // @[Conditional.scala 39:67]
  wire  _GEN_1542 = _T_83 ? valid_0_0 : _GEN_1470; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1543 = _T_83 ? valid_0_1 : _GEN_1471; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1544 = _T_83 ? valid_0_2 : _GEN_1472; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1545 = _T_83 ? valid_0_3 : _GEN_1473; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1546 = _T_83 ? valid_0_4 : _GEN_1474; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1547 = _T_83 ? valid_0_5 : _GEN_1475; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1548 = _T_83 ? valid_0_6 : _GEN_1476; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1549 = _T_83 ? valid_0_7 : _GEN_1477; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1550 = _T_83 ? valid_0_8 : _GEN_1478; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1551 = _T_83 ? valid_0_9 : _GEN_1479; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1552 = _T_83 ? valid_0_10 : _GEN_1480; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1553 = _T_83 ? valid_0_11 : _GEN_1481; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1554 = _T_83 ? valid_0_12 : _GEN_1482; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1555 = _T_83 ? valid_0_13 : _GEN_1483; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1556 = _T_83 ? valid_0_14 : _GEN_1484; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1557 = _T_83 ? valid_0_15 : _GEN_1485; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1558 = _T_83 ? valid_1_0 : _GEN_1486; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1559 = _T_83 ? valid_1_1 : _GEN_1487; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1560 = _T_83 ? valid_1_2 : _GEN_1488; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1561 = _T_83 ? valid_1_3 : _GEN_1489; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1562 = _T_83 ? valid_1_4 : _GEN_1490; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1563 = _T_83 ? valid_1_5 : _GEN_1491; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1564 = _T_83 ? valid_1_6 : _GEN_1492; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1565 = _T_83 ? valid_1_7 : _GEN_1493; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1566 = _T_83 ? valid_1_8 : _GEN_1494; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1567 = _T_83 ? valid_1_9 : _GEN_1495; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1568 = _T_83 ? valid_1_10 : _GEN_1496; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1569 = _T_83 ? valid_1_11 : _GEN_1497; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1570 = _T_83 ? valid_1_12 : _GEN_1498; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1571 = _T_83 ? valid_1_13 : _GEN_1499; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1572 = _T_83 ? valid_1_14 : _GEN_1500; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1573 = _T_83 ? valid_1_15 : _GEN_1501; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1574 = _T_83 ? valid_2_0 : _GEN_1502; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1575 = _T_83 ? valid_2_1 : _GEN_1503; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1576 = _T_83 ? valid_2_2 : _GEN_1504; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1577 = _T_83 ? valid_2_3 : _GEN_1505; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1578 = _T_83 ? valid_2_4 : _GEN_1506; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1579 = _T_83 ? valid_2_5 : _GEN_1507; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1580 = _T_83 ? valid_2_6 : _GEN_1508; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1581 = _T_83 ? valid_2_7 : _GEN_1509; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1582 = _T_83 ? valid_2_8 : _GEN_1510; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1583 = _T_83 ? valid_2_9 : _GEN_1511; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1584 = _T_83 ? valid_2_10 : _GEN_1512; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1585 = _T_83 ? valid_2_11 : _GEN_1513; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1586 = _T_83 ? valid_2_12 : _GEN_1514; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1587 = _T_83 ? valid_2_13 : _GEN_1515; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1588 = _T_83 ? valid_2_14 : _GEN_1516; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1589 = _T_83 ? valid_2_15 : _GEN_1517; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1590 = _T_83 ? valid_3_0 : _GEN_1518; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1591 = _T_83 ? valid_3_1 : _GEN_1519; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1592 = _T_83 ? valid_3_2 : _GEN_1520; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1593 = _T_83 ? valid_3_3 : _GEN_1521; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1594 = _T_83 ? valid_3_4 : _GEN_1522; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1595 = _T_83 ? valid_3_5 : _GEN_1523; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1596 = _T_83 ? valid_3_6 : _GEN_1524; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1597 = _T_83 ? valid_3_7 : _GEN_1525; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1598 = _T_83 ? valid_3_8 : _GEN_1526; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1599 = _T_83 ? valid_3_9 : _GEN_1527; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1600 = _T_83 ? valid_3_10 : _GEN_1528; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1601 = _T_83 ? valid_3_11 : _GEN_1529; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1602 = _T_83 ? valid_3_12 : _GEN_1530; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1603 = _T_83 ? valid_3_13 : _GEN_1531; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1604 = _T_83 ? valid_3_14 : _GEN_1532; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1605 = _T_83 ? valid_3_15 : _GEN_1533; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1606 = _T_83 ? axiWaddrEn : _GEN_1534; // @[Conditional.scala 39:67 dcache.scala 221:34]
  wire [1:0] _GEN_1607 = _T_83 ? _GEN_129 : _GEN_1535; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_1608 = _T_83 ? _GEN_133 : _GEN_1536; // @[Conditional.scala 39:67]
  wire  _GEN_1609 = _T_81 ? _GEN_1269 : axiWdataEn; // @[Conditional.scala 39:67 dcache.scala 224:34]
  wire [2:0] _GEN_1610 = _T_81 ? _GEN_1268 : offset; // @[Conditional.scala 39:67 dcache.scala 111:34]
  wire [2:0] _GEN_1611 = _T_81 ? _GEN_1270 : _GEN_1540; // @[Conditional.scala 39:67]
  wire  _GEN_1612 = _T_81 ? _GEN_1271 : _GEN_1542; // @[Conditional.scala 39:67]
  wire  _GEN_1613 = _T_81 ? _GEN_1272 : _GEN_1543; // @[Conditional.scala 39:67]
  wire  _GEN_1614 = _T_81 ? _GEN_1273 : _GEN_1544; // @[Conditional.scala 39:67]
  wire  _GEN_1615 = _T_81 ? _GEN_1274 : _GEN_1545; // @[Conditional.scala 39:67]
  wire  _GEN_1616 = _T_81 ? _GEN_1275 : _GEN_1546; // @[Conditional.scala 39:67]
  wire  _GEN_1617 = _T_81 ? _GEN_1276 : _GEN_1547; // @[Conditional.scala 39:67]
  wire  _GEN_1618 = _T_81 ? _GEN_1277 : _GEN_1548; // @[Conditional.scala 39:67]
  wire  _GEN_1619 = _T_81 ? _GEN_1278 : _GEN_1549; // @[Conditional.scala 39:67]
  wire  _GEN_1620 = _T_81 ? _GEN_1279 : _GEN_1550; // @[Conditional.scala 39:67]
  wire  _GEN_1621 = _T_81 ? _GEN_1280 : _GEN_1551; // @[Conditional.scala 39:67]
  wire  _GEN_1622 = _T_81 ? _GEN_1281 : _GEN_1552; // @[Conditional.scala 39:67]
  wire  _GEN_1623 = _T_81 ? _GEN_1282 : _GEN_1553; // @[Conditional.scala 39:67]
  wire  _GEN_1624 = _T_81 ? _GEN_1283 : _GEN_1554; // @[Conditional.scala 39:67]
  wire  _GEN_1625 = _T_81 ? _GEN_1284 : _GEN_1555; // @[Conditional.scala 39:67]
  wire  _GEN_1626 = _T_81 ? _GEN_1285 : _GEN_1556; // @[Conditional.scala 39:67]
  wire  _GEN_1627 = _T_81 ? _GEN_1286 : _GEN_1557; // @[Conditional.scala 39:67]
  wire  _GEN_1628 = _T_81 ? _GEN_1287 : _GEN_1558; // @[Conditional.scala 39:67]
  wire  _GEN_1629 = _T_81 ? _GEN_1288 : _GEN_1559; // @[Conditional.scala 39:67]
  wire  _GEN_1630 = _T_81 ? _GEN_1289 : _GEN_1560; // @[Conditional.scala 39:67]
  wire  _GEN_1631 = _T_81 ? _GEN_1290 : _GEN_1561; // @[Conditional.scala 39:67]
  wire  _GEN_1632 = _T_81 ? _GEN_1291 : _GEN_1562; // @[Conditional.scala 39:67]
  wire  _GEN_1633 = _T_81 ? _GEN_1292 : _GEN_1563; // @[Conditional.scala 39:67]
  wire  _GEN_1634 = _T_81 ? _GEN_1293 : _GEN_1564; // @[Conditional.scala 39:67]
  wire  _GEN_1635 = _T_81 ? _GEN_1294 : _GEN_1565; // @[Conditional.scala 39:67]
  wire  _GEN_1636 = _T_81 ? _GEN_1295 : _GEN_1566; // @[Conditional.scala 39:67]
  wire  _GEN_1637 = _T_81 ? _GEN_1296 : _GEN_1567; // @[Conditional.scala 39:67]
  wire  _GEN_1638 = _T_81 ? _GEN_1297 : _GEN_1568; // @[Conditional.scala 39:67]
  wire  _GEN_1639 = _T_81 ? _GEN_1298 : _GEN_1569; // @[Conditional.scala 39:67]
  wire  _GEN_1640 = _T_81 ? _GEN_1299 : _GEN_1570; // @[Conditional.scala 39:67]
  wire  _GEN_1641 = _T_81 ? _GEN_1300 : _GEN_1571; // @[Conditional.scala 39:67]
  wire  _GEN_1642 = _T_81 ? _GEN_1301 : _GEN_1572; // @[Conditional.scala 39:67]
  wire  _GEN_1643 = _T_81 ? _GEN_1302 : _GEN_1573; // @[Conditional.scala 39:67]
  wire  _GEN_1644 = _T_81 ? _GEN_1303 : _GEN_1574; // @[Conditional.scala 39:67]
  wire  _GEN_1645 = _T_81 ? _GEN_1304 : _GEN_1575; // @[Conditional.scala 39:67]
  wire  _GEN_1646 = _T_81 ? _GEN_1305 : _GEN_1576; // @[Conditional.scala 39:67]
  wire  _GEN_1647 = _T_81 ? _GEN_1306 : _GEN_1577; // @[Conditional.scala 39:67]
  wire  _GEN_1648 = _T_81 ? _GEN_1307 : _GEN_1578; // @[Conditional.scala 39:67]
  wire  _GEN_1649 = _T_81 ? _GEN_1308 : _GEN_1579; // @[Conditional.scala 39:67]
  wire  _GEN_1650 = _T_81 ? _GEN_1309 : _GEN_1580; // @[Conditional.scala 39:67]
  wire  _GEN_1651 = _T_81 ? _GEN_1310 : _GEN_1581; // @[Conditional.scala 39:67]
  wire  _GEN_1652 = _T_81 ? _GEN_1311 : _GEN_1582; // @[Conditional.scala 39:67]
  wire  _GEN_1653 = _T_81 ? _GEN_1312 : _GEN_1583; // @[Conditional.scala 39:67]
  wire  _GEN_1654 = _T_81 ? _GEN_1313 : _GEN_1584; // @[Conditional.scala 39:67]
  wire  _GEN_1655 = _T_81 ? _GEN_1314 : _GEN_1585; // @[Conditional.scala 39:67]
  wire  _GEN_1656 = _T_81 ? _GEN_1315 : _GEN_1586; // @[Conditional.scala 39:67]
  wire  _GEN_1657 = _T_81 ? _GEN_1316 : _GEN_1587; // @[Conditional.scala 39:67]
  wire  _GEN_1658 = _T_81 ? _GEN_1317 : _GEN_1588; // @[Conditional.scala 39:67]
  wire  _GEN_1659 = _T_81 ? _GEN_1318 : _GEN_1589; // @[Conditional.scala 39:67]
  wire  _GEN_1660 = _T_81 ? _GEN_1319 : _GEN_1590; // @[Conditional.scala 39:67]
  wire  _GEN_1661 = _T_81 ? _GEN_1320 : _GEN_1591; // @[Conditional.scala 39:67]
  wire  _GEN_1662 = _T_81 ? _GEN_1321 : _GEN_1592; // @[Conditional.scala 39:67]
  wire  _GEN_1663 = _T_81 ? _GEN_1322 : _GEN_1593; // @[Conditional.scala 39:67]
  wire  _GEN_1664 = _T_81 ? _GEN_1323 : _GEN_1594; // @[Conditional.scala 39:67]
  wire  _GEN_1665 = _T_81 ? _GEN_1324 : _GEN_1595; // @[Conditional.scala 39:67]
  wire  _GEN_1666 = _T_81 ? _GEN_1325 : _GEN_1596; // @[Conditional.scala 39:67]
  wire  _GEN_1667 = _T_81 ? _GEN_1326 : _GEN_1597; // @[Conditional.scala 39:67]
  wire  _GEN_1668 = _T_81 ? _GEN_1327 : _GEN_1598; // @[Conditional.scala 39:67]
  wire  _GEN_1669 = _T_81 ? _GEN_1328 : _GEN_1599; // @[Conditional.scala 39:67]
  wire  _GEN_1670 = _T_81 ? _GEN_1329 : _GEN_1600; // @[Conditional.scala 39:67]
  wire  _GEN_1671 = _T_81 ? _GEN_1330 : _GEN_1601; // @[Conditional.scala 39:67]
  wire  _GEN_1672 = _T_81 ? _GEN_1331 : _GEN_1602; // @[Conditional.scala 39:67]
  wire  _GEN_1673 = _T_81 ? _GEN_1332 : _GEN_1603; // @[Conditional.scala 39:67]
  wire  _GEN_1674 = _T_81 ? _GEN_1333 : _GEN_1604; // @[Conditional.scala 39:67]
  wire  _GEN_1675 = _T_81 ? _GEN_1334 : _GEN_1605; // @[Conditional.scala 39:67]
  wire  _GEN_1676 = _T_81 ? _GEN_1335 : _GEN_390; // @[Conditional.scala 39:67]
  wire  _GEN_1677 = _T_81 ? _GEN_1336 : _GEN_391; // @[Conditional.scala 39:67]
  wire  _GEN_1678 = _T_81 ? _GEN_1337 : _GEN_392; // @[Conditional.scala 39:67]
  wire  _GEN_1679 = _T_81 ? _GEN_1338 : _GEN_393; // @[Conditional.scala 39:67]
  wire  _GEN_1680 = _T_81 ? _GEN_1339 : _GEN_394; // @[Conditional.scala 39:67]
  wire  _GEN_1681 = _T_81 ? _GEN_1340 : _GEN_395; // @[Conditional.scala 39:67]
  wire  _GEN_1682 = _T_81 ? _GEN_1341 : _GEN_396; // @[Conditional.scala 39:67]
  wire  _GEN_1683 = _T_81 ? _GEN_1342 : _GEN_397; // @[Conditional.scala 39:67]
  wire  _GEN_1684 = _T_81 ? _GEN_1343 : _GEN_398; // @[Conditional.scala 39:67]
  wire  _GEN_1685 = _T_81 ? _GEN_1344 : _GEN_399; // @[Conditional.scala 39:67]
  wire  _GEN_1686 = _T_81 ? _GEN_1345 : _GEN_400; // @[Conditional.scala 39:67]
  wire  _GEN_1687 = _T_81 ? _GEN_1346 : _GEN_401; // @[Conditional.scala 39:67]
  wire  _GEN_1688 = _T_81 ? _GEN_1347 : _GEN_402; // @[Conditional.scala 39:67]
  wire  _GEN_1689 = _T_81 ? _GEN_1348 : _GEN_403; // @[Conditional.scala 39:67]
  wire  _GEN_1690 = _T_81 ? _GEN_1349 : _GEN_404; // @[Conditional.scala 39:67]
  wire  _GEN_1691 = _T_81 ? _GEN_1350 : _GEN_405; // @[Conditional.scala 39:67]
  wire  _GEN_1692 = _T_81 ? _GEN_1351 : _GEN_406; // @[Conditional.scala 39:67]
  wire  _GEN_1693 = _T_81 ? _GEN_1352 : _GEN_407; // @[Conditional.scala 39:67]
  wire  _GEN_1694 = _T_81 ? _GEN_1353 : _GEN_408; // @[Conditional.scala 39:67]
  wire  _GEN_1695 = _T_81 ? _GEN_1354 : _GEN_409; // @[Conditional.scala 39:67]
  wire  _GEN_1696 = _T_81 ? _GEN_1355 : _GEN_410; // @[Conditional.scala 39:67]
  wire  _GEN_1697 = _T_81 ? _GEN_1356 : _GEN_411; // @[Conditional.scala 39:67]
  wire  _GEN_1698 = _T_81 ? _GEN_1357 : _GEN_412; // @[Conditional.scala 39:67]
  wire  _GEN_1699 = _T_81 ? _GEN_1358 : _GEN_413; // @[Conditional.scala 39:67]
  wire  _GEN_1700 = _T_81 ? _GEN_1359 : _GEN_414; // @[Conditional.scala 39:67]
  wire  _GEN_1701 = _T_81 ? _GEN_1360 : _GEN_415; // @[Conditional.scala 39:67]
  wire  _GEN_1702 = _T_81 ? _GEN_1361 : _GEN_416; // @[Conditional.scala 39:67]
  wire  _GEN_1703 = _T_81 ? _GEN_1362 : _GEN_417; // @[Conditional.scala 39:67]
  wire  _GEN_1704 = _T_81 ? _GEN_1363 : _GEN_418; // @[Conditional.scala 39:67]
  wire  _GEN_1705 = _T_81 ? _GEN_1364 : _GEN_419; // @[Conditional.scala 39:67]
  wire  _GEN_1706 = _T_81 ? _GEN_1365 : _GEN_420; // @[Conditional.scala 39:67]
  wire  _GEN_1707 = _T_81 ? _GEN_1366 : _GEN_421; // @[Conditional.scala 39:67]
  wire  _GEN_1708 = _T_81 ? _GEN_1367 : _GEN_422; // @[Conditional.scala 39:67]
  wire  _GEN_1709 = _T_81 ? _GEN_1368 : _GEN_423; // @[Conditional.scala 39:67]
  wire  _GEN_1710 = _T_81 ? _GEN_1369 : _GEN_424; // @[Conditional.scala 39:67]
  wire  _GEN_1711 = _T_81 ? _GEN_1370 : _GEN_425; // @[Conditional.scala 39:67]
  wire  _GEN_1712 = _T_81 ? _GEN_1371 : _GEN_426; // @[Conditional.scala 39:67]
  wire  _GEN_1713 = _T_81 ? _GEN_1372 : _GEN_427; // @[Conditional.scala 39:67]
  wire  _GEN_1714 = _T_81 ? _GEN_1373 : _GEN_428; // @[Conditional.scala 39:67]
  wire  _GEN_1715 = _T_81 ? _GEN_1374 : _GEN_429; // @[Conditional.scala 39:67]
  wire  _GEN_1716 = _T_81 ? _GEN_1375 : _GEN_430; // @[Conditional.scala 39:67]
  wire  _GEN_1717 = _T_81 ? _GEN_1376 : _GEN_431; // @[Conditional.scala 39:67]
  wire  _GEN_1718 = _T_81 ? _GEN_1377 : _GEN_432; // @[Conditional.scala 39:67]
  wire  _GEN_1719 = _T_81 ? _GEN_1378 : _GEN_433; // @[Conditional.scala 39:67]
  wire  _GEN_1720 = _T_81 ? _GEN_1379 : _GEN_434; // @[Conditional.scala 39:67]
  wire  _GEN_1721 = _T_81 ? _GEN_1380 : _GEN_435; // @[Conditional.scala 39:67]
  wire  _GEN_1722 = _T_81 ? _GEN_1381 : _GEN_436; // @[Conditional.scala 39:67]
  wire  _GEN_1723 = _T_81 ? _GEN_1382 : _GEN_437; // @[Conditional.scala 39:67]
  wire  _GEN_1724 = _T_81 ? _GEN_1383 : _GEN_438; // @[Conditional.scala 39:67]
  wire  _GEN_1725 = _T_81 ? _GEN_1384 : _GEN_439; // @[Conditional.scala 39:67]
  wire  _GEN_1726 = _T_81 ? _GEN_1385 : _GEN_440; // @[Conditional.scala 39:67]
  wire  _GEN_1727 = _T_81 ? _GEN_1386 : _GEN_441; // @[Conditional.scala 39:67]
  wire  _GEN_1728 = _T_81 ? _GEN_1387 : _GEN_442; // @[Conditional.scala 39:67]
  wire  _GEN_1729 = _T_81 ? _GEN_1388 : _GEN_443; // @[Conditional.scala 39:67]
  wire  _GEN_1730 = _T_81 ? _GEN_1389 : _GEN_444; // @[Conditional.scala 39:67]
  wire  _GEN_1731 = _T_81 ? _GEN_1390 : _GEN_445; // @[Conditional.scala 39:67]
  wire  _GEN_1732 = _T_81 ? _GEN_1391 : _GEN_446; // @[Conditional.scala 39:67]
  wire  _GEN_1733 = _T_81 ? _GEN_1392 : _GEN_447; // @[Conditional.scala 39:67]
  wire  _GEN_1734 = _T_81 ? _GEN_1393 : _GEN_448; // @[Conditional.scala 39:67]
  wire  _GEN_1735 = _T_81 ? _GEN_1394 : _GEN_449; // @[Conditional.scala 39:67]
  wire  _GEN_1736 = _T_81 ? _GEN_1395 : _GEN_450; // @[Conditional.scala 39:67]
  wire  _GEN_1737 = _T_81 ? _GEN_1396 : _GEN_451; // @[Conditional.scala 39:67]
  wire  _GEN_1738 = _T_81 ? _GEN_1397 : _GEN_452; // @[Conditional.scala 39:67]
  wire  _GEN_1739 = _T_81 ? _GEN_1398 : _GEN_453; // @[Conditional.scala 39:67]
  wire  _GEN_1742 = _T_81 ? wait_r : _GEN_1539; // @[Conditional.scala 39:67 dcache.scala 96:30]
  wire  _GEN_1743 = _T_81 ? _GEN_134 : _GEN_1541; // @[Conditional.scala 39:67]
  wire  _GEN_1744 = _T_81 ? axiWaddrEn : _GEN_1606; // @[Conditional.scala 39:67 dcache.scala 221:34]
  wire [1:0] _GEN_1745 = _T_81 ? _GEN_129 : _GEN_1607; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_1746 = _T_81 ? _GEN_133 : _GEN_1608; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_1747 = _T_79 ? 3'h0 : _GEN_1610; // @[Conditional.scala 39:67 dcache.scala 281:20]
  wire [2:0] _GEN_1748 = _T_79 ? _GEN_1007 : _GEN_1611; // @[Conditional.scala 39:67]
  wire  _GEN_1749 = _T_79 ? _GEN_1008 : _GEN_1744; // @[Conditional.scala 39:67]
  wire  _GEN_1750 = _T_79 ? _GEN_1009 : _GEN_1609; // @[Conditional.scala 39:67]
  wire  _GEN_1751 = _T_79 ? valid_0_0 : _GEN_1612; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1752 = _T_79 ? valid_0_1 : _GEN_1613; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1753 = _T_79 ? valid_0_2 : _GEN_1614; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1754 = _T_79 ? valid_0_3 : _GEN_1615; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1755 = _T_79 ? valid_0_4 : _GEN_1616; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1756 = _T_79 ? valid_0_5 : _GEN_1617; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1757 = _T_79 ? valid_0_6 : _GEN_1618; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1758 = _T_79 ? valid_0_7 : _GEN_1619; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1759 = _T_79 ? valid_0_8 : _GEN_1620; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1760 = _T_79 ? valid_0_9 : _GEN_1621; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1761 = _T_79 ? valid_0_10 : _GEN_1622; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1762 = _T_79 ? valid_0_11 : _GEN_1623; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1763 = _T_79 ? valid_0_12 : _GEN_1624; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1764 = _T_79 ? valid_0_13 : _GEN_1625; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1765 = _T_79 ? valid_0_14 : _GEN_1626; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1766 = _T_79 ? valid_0_15 : _GEN_1627; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1767 = _T_79 ? valid_1_0 : _GEN_1628; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1768 = _T_79 ? valid_1_1 : _GEN_1629; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1769 = _T_79 ? valid_1_2 : _GEN_1630; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1770 = _T_79 ? valid_1_3 : _GEN_1631; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1771 = _T_79 ? valid_1_4 : _GEN_1632; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1772 = _T_79 ? valid_1_5 : _GEN_1633; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1773 = _T_79 ? valid_1_6 : _GEN_1634; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1774 = _T_79 ? valid_1_7 : _GEN_1635; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1775 = _T_79 ? valid_1_8 : _GEN_1636; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1776 = _T_79 ? valid_1_9 : _GEN_1637; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1777 = _T_79 ? valid_1_10 : _GEN_1638; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1778 = _T_79 ? valid_1_11 : _GEN_1639; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1779 = _T_79 ? valid_1_12 : _GEN_1640; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1780 = _T_79 ? valid_1_13 : _GEN_1641; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1781 = _T_79 ? valid_1_14 : _GEN_1642; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1782 = _T_79 ? valid_1_15 : _GEN_1643; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1783 = _T_79 ? valid_2_0 : _GEN_1644; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1784 = _T_79 ? valid_2_1 : _GEN_1645; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1785 = _T_79 ? valid_2_2 : _GEN_1646; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1786 = _T_79 ? valid_2_3 : _GEN_1647; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1787 = _T_79 ? valid_2_4 : _GEN_1648; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1788 = _T_79 ? valid_2_5 : _GEN_1649; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1789 = _T_79 ? valid_2_6 : _GEN_1650; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1790 = _T_79 ? valid_2_7 : _GEN_1651; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1791 = _T_79 ? valid_2_8 : _GEN_1652; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1792 = _T_79 ? valid_2_9 : _GEN_1653; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1793 = _T_79 ? valid_2_10 : _GEN_1654; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1794 = _T_79 ? valid_2_11 : _GEN_1655; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1795 = _T_79 ? valid_2_12 : _GEN_1656; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1796 = _T_79 ? valid_2_13 : _GEN_1657; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1797 = _T_79 ? valid_2_14 : _GEN_1658; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1798 = _T_79 ? valid_2_15 : _GEN_1659; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1799 = _T_79 ? valid_3_0 : _GEN_1660; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1800 = _T_79 ? valid_3_1 : _GEN_1661; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1801 = _T_79 ? valid_3_2 : _GEN_1662; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1802 = _T_79 ? valid_3_3 : _GEN_1663; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1803 = _T_79 ? valid_3_4 : _GEN_1664; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1804 = _T_79 ? valid_3_5 : _GEN_1665; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1805 = _T_79 ? valid_3_6 : _GEN_1666; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1806 = _T_79 ? valid_3_7 : _GEN_1667; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1807 = _T_79 ? valid_3_8 : _GEN_1668; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1808 = _T_79 ? valid_3_9 : _GEN_1669; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1809 = _T_79 ? valid_3_10 : _GEN_1670; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1810 = _T_79 ? valid_3_11 : _GEN_1671; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1811 = _T_79 ? valid_3_12 : _GEN_1672; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1812 = _T_79 ? valid_3_13 : _GEN_1673; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1813 = _T_79 ? valid_3_14 : _GEN_1674; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1814 = _T_79 ? valid_3_15 : _GEN_1675; // @[Conditional.scala 39:67 dcache.scala 93:26]
  wire  _GEN_1815 = _T_79 ? _GEN_390 : _GEN_1676; // @[Conditional.scala 39:67]
  wire  _GEN_1816 = _T_79 ? _GEN_391 : _GEN_1677; // @[Conditional.scala 39:67]
  wire  _GEN_1817 = _T_79 ? _GEN_392 : _GEN_1678; // @[Conditional.scala 39:67]
  wire  _GEN_1818 = _T_79 ? _GEN_393 : _GEN_1679; // @[Conditional.scala 39:67]
  wire  _GEN_1819 = _T_79 ? _GEN_394 : _GEN_1680; // @[Conditional.scala 39:67]
  wire  _GEN_1820 = _T_79 ? _GEN_395 : _GEN_1681; // @[Conditional.scala 39:67]
  wire  _GEN_1821 = _T_79 ? _GEN_396 : _GEN_1682; // @[Conditional.scala 39:67]
  wire  _GEN_1822 = _T_79 ? _GEN_397 : _GEN_1683; // @[Conditional.scala 39:67]
  wire  _GEN_1823 = _T_79 ? _GEN_398 : _GEN_1684; // @[Conditional.scala 39:67]
  wire  _GEN_1824 = _T_79 ? _GEN_399 : _GEN_1685; // @[Conditional.scala 39:67]
  wire  _GEN_1825 = _T_79 ? _GEN_400 : _GEN_1686; // @[Conditional.scala 39:67]
  wire  _GEN_1826 = _T_79 ? _GEN_401 : _GEN_1687; // @[Conditional.scala 39:67]
  wire  _GEN_1827 = _T_79 ? _GEN_402 : _GEN_1688; // @[Conditional.scala 39:67]
  wire  _GEN_1828 = _T_79 ? _GEN_403 : _GEN_1689; // @[Conditional.scala 39:67]
  wire  _GEN_1829 = _T_79 ? _GEN_404 : _GEN_1690; // @[Conditional.scala 39:67]
  wire  _GEN_1830 = _T_79 ? _GEN_405 : _GEN_1691; // @[Conditional.scala 39:67]
  wire  _GEN_1831 = _T_79 ? _GEN_406 : _GEN_1692; // @[Conditional.scala 39:67]
  wire  _GEN_1832 = _T_79 ? _GEN_407 : _GEN_1693; // @[Conditional.scala 39:67]
  wire  _GEN_1833 = _T_79 ? _GEN_408 : _GEN_1694; // @[Conditional.scala 39:67]
  wire  _GEN_1834 = _T_79 ? _GEN_409 : _GEN_1695; // @[Conditional.scala 39:67]
  wire  _GEN_1835 = _T_79 ? _GEN_410 : _GEN_1696; // @[Conditional.scala 39:67]
  wire  _GEN_1836 = _T_79 ? _GEN_411 : _GEN_1697; // @[Conditional.scala 39:67]
  wire  _GEN_1837 = _T_79 ? _GEN_412 : _GEN_1698; // @[Conditional.scala 39:67]
  wire  _GEN_1838 = _T_79 ? _GEN_413 : _GEN_1699; // @[Conditional.scala 39:67]
  wire  _GEN_1839 = _T_79 ? _GEN_414 : _GEN_1700; // @[Conditional.scala 39:67]
  wire  _GEN_1840 = _T_79 ? _GEN_415 : _GEN_1701; // @[Conditional.scala 39:67]
  wire  _GEN_1841 = _T_79 ? _GEN_416 : _GEN_1702; // @[Conditional.scala 39:67]
  wire  _GEN_1842 = _T_79 ? _GEN_417 : _GEN_1703; // @[Conditional.scala 39:67]
  wire  _GEN_1843 = _T_79 ? _GEN_418 : _GEN_1704; // @[Conditional.scala 39:67]
  wire  _GEN_1844 = _T_79 ? _GEN_419 : _GEN_1705; // @[Conditional.scala 39:67]
  wire  _GEN_1845 = _T_79 ? _GEN_420 : _GEN_1706; // @[Conditional.scala 39:67]
  wire  _GEN_1846 = _T_79 ? _GEN_421 : _GEN_1707; // @[Conditional.scala 39:67]
  wire  _GEN_1847 = _T_79 ? _GEN_422 : _GEN_1708; // @[Conditional.scala 39:67]
  wire  _GEN_1848 = _T_79 ? _GEN_423 : _GEN_1709; // @[Conditional.scala 39:67]
  wire  _GEN_1849 = _T_79 ? _GEN_424 : _GEN_1710; // @[Conditional.scala 39:67]
  wire  _GEN_1850 = _T_79 ? _GEN_425 : _GEN_1711; // @[Conditional.scala 39:67]
  wire  _GEN_1851 = _T_79 ? _GEN_426 : _GEN_1712; // @[Conditional.scala 39:67]
  wire  _GEN_1852 = _T_79 ? _GEN_427 : _GEN_1713; // @[Conditional.scala 39:67]
  wire  _GEN_1853 = _T_79 ? _GEN_428 : _GEN_1714; // @[Conditional.scala 39:67]
  wire  _GEN_1854 = _T_79 ? _GEN_429 : _GEN_1715; // @[Conditional.scala 39:67]
  wire  _GEN_1855 = _T_79 ? _GEN_430 : _GEN_1716; // @[Conditional.scala 39:67]
  wire  _GEN_1856 = _T_79 ? _GEN_431 : _GEN_1717; // @[Conditional.scala 39:67]
  wire  _GEN_1857 = _T_79 ? _GEN_432 : _GEN_1718; // @[Conditional.scala 39:67]
  wire  _GEN_1858 = _T_79 ? _GEN_433 : _GEN_1719; // @[Conditional.scala 39:67]
  wire  _GEN_1859 = _T_79 ? _GEN_434 : _GEN_1720; // @[Conditional.scala 39:67]
  wire  _GEN_1860 = _T_79 ? _GEN_435 : _GEN_1721; // @[Conditional.scala 39:67]
  wire  _GEN_1861 = _T_79 ? _GEN_436 : _GEN_1722; // @[Conditional.scala 39:67]
  wire  _GEN_1862 = _T_79 ? _GEN_437 : _GEN_1723; // @[Conditional.scala 39:67]
  wire  _GEN_1863 = _T_79 ? _GEN_438 : _GEN_1724; // @[Conditional.scala 39:67]
  wire  _GEN_1864 = _T_79 ? _GEN_439 : _GEN_1725; // @[Conditional.scala 39:67]
  wire  _GEN_1865 = _T_79 ? _GEN_440 : _GEN_1726; // @[Conditional.scala 39:67]
  wire  _GEN_1866 = _T_79 ? _GEN_441 : _GEN_1727; // @[Conditional.scala 39:67]
  wire  _GEN_1867 = _T_79 ? _GEN_442 : _GEN_1728; // @[Conditional.scala 39:67]
  wire  _GEN_1868 = _T_79 ? _GEN_443 : _GEN_1729; // @[Conditional.scala 39:67]
  wire  _GEN_1869 = _T_79 ? _GEN_444 : _GEN_1730; // @[Conditional.scala 39:67]
  wire  _GEN_1870 = _T_79 ? _GEN_445 : _GEN_1731; // @[Conditional.scala 39:67]
  wire  _GEN_1871 = _T_79 ? _GEN_446 : _GEN_1732; // @[Conditional.scala 39:67]
  wire  _GEN_1872 = _T_79 ? _GEN_447 : _GEN_1733; // @[Conditional.scala 39:67]
  wire  _GEN_1873 = _T_79 ? _GEN_448 : _GEN_1734; // @[Conditional.scala 39:67]
  wire  _GEN_1874 = _T_79 ? _GEN_449 : _GEN_1735; // @[Conditional.scala 39:67]
  wire  _GEN_1875 = _T_79 ? _GEN_450 : _GEN_1736; // @[Conditional.scala 39:67]
  wire  _GEN_1876 = _T_79 ? _GEN_451 : _GEN_1737; // @[Conditional.scala 39:67]
  wire  _GEN_1877 = _T_79 ? _GEN_452 : _GEN_1738; // @[Conditional.scala 39:67]
  wire  _GEN_1878 = _T_79 ? _GEN_453 : _GEN_1739; // @[Conditional.scala 39:67]
  wire  _GEN_1881 = _T_79 ? wait_r : _GEN_1742; // @[Conditional.scala 39:67 dcache.scala 96:30]
  wire  _GEN_1882 = _T_79 ? _GEN_134 : _GEN_1743; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_1883 = _T_79 ? _GEN_129 : _GEN_1745; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_1884 = _T_79 ? _GEN_133 : _GEN_1746; // @[Conditional.scala 39:67]
  wire  _GEN_2295 = _T_68 & _GEN_605; // @[Conditional.scala 40:58 dcache.scala 102:13]
  ysyx_210539_MaxPeriodFibonacciLFSR matchWay_prng ( // @[PRNG.scala 82:22]
    .clock(matchWay_prng_clock),
    .reset(matchWay_prng_reset),
    .io_out_0(matchWay_prng_io_out_0),
    .io_out_1(matchWay_prng_io_out_1),
    .io_out_2(matchWay_prng_io_out_2)
  );
  assign io_dataAxi_wa_valid = axiWaddrEn; // @[dcache.scala 330:30]
  assign io_dataAxi_wa_bits_addr = {axiWaddr_hi,6'h0}; // @[Cat.scala 30:58]
  assign io_dataAxi_wd_valid = axiWdataEn; // @[dcache.scala 336:30]
  assign io_dataAxi_wd_bits_data = offset[0] ? rdata128[127:64] : rdata128[63:0]; // @[dcache.scala 223:30]
  assign io_dataAxi_wd_bits_last = offset == 3'h7; // @[dcache.scala 225:34]
  assign io_dataAxi_ra_valid = axiRaddrEn; // @[dcache.scala 322:30]
  assign io_dataAxi_ra_bits_addr = cur_addr & 32'hffffffc0; // @[dcache.scala 219:36]
  assign io_dcRW_rdata = _io_dcRW_rdata_T_32[63:0]; // @[dcache.scala 161:19]
  assign io_dcRW_rvalid = valid_r; // @[dcache.scala 106:20]
  assign io_dcRW_ready = valid_in & ~wait_r; // @[dcache.scala 105:31]
  assign io_flush_out = flush_r; // @[dcache.scala 107:18]
  assign io_dc2sr0_addr = state == 3'h0 | state == 3'h5 ? cur_ram_addr : cur_axi_addr; // @[dcache.scala 190:26]
  assign io_dc2sr0_cen = ~(_GEN_129 == 2'h0 & (wait_r | hs_in | flush_r)); // @[dcache.scala 194:22]
  assign io_dc2sr0_wen = ~wen; // @[dcache.scala 198:22]
  assign io_dc2sr0_wmask = ~mask; // @[dcache.scala 207:24]
  assign io_dc2sr0_wdata = _io_dc2sr0_wdata_T_4[127:0]; // @[dcache.scala 202:21]
  assign io_dc2sr1_addr = io_dc2sr0_addr; // @[dcache.scala 191:20]
  assign io_dc2sr1_cen = ~(_GEN_129 == 2'h1 & _io_dc2sr0_cen_T_2); // @[dcache.scala 195:22]
  assign io_dc2sr1_wen = io_dc2sr0_wen; // @[dcache.scala 199:19]
  assign io_dc2sr1_wmask = io_dc2sr0_wmask; // @[dcache.scala 208:21]
  assign io_dc2sr1_wdata = io_dc2sr0_wdata; // @[dcache.scala 204:21]
  assign io_dc2sr2_addr = io_dc2sr0_addr; // @[dcache.scala 192:20]
  assign io_dc2sr2_cen = ~(_GEN_129 == 2'h2 & _io_dc2sr0_cen_T_2); // @[dcache.scala 196:22]
  assign io_dc2sr2_wen = io_dc2sr0_wen; // @[dcache.scala 200:19]
  assign io_dc2sr2_wmask = io_dc2sr0_wmask; // @[dcache.scala 209:21]
  assign io_dc2sr2_wdata = io_dc2sr0_wdata; // @[dcache.scala 205:21]
  assign io_dc2sr3_addr = io_dc2sr0_addr; // @[dcache.scala 193:20]
  assign io_dc2sr3_cen = ~(_GEN_129 == 2'h3 & _io_dc2sr0_cen_T_2); // @[dcache.scala 197:22]
  assign io_dc2sr3_wen = io_dc2sr0_wen; // @[dcache.scala 201:19]
  assign io_dc2sr3_wmask = io_dc2sr0_wmask; // @[dcache.scala 210:21]
  assign io_dc2sr3_wdata = io_dc2sr0_wdata; // @[dcache.scala 206:21]
  assign matchWay_prng_clock = clock;
  assign matchWay_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[dcache.scala 92:26]
      tag_0_0 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_0_0 <= _GEN_878;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_0_1 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_0_1 <= _GEN_879;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_0_2 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_0_2 <= _GEN_880;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_0_3 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_0_3 <= _GEN_881;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_0_4 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_0_4 <= _GEN_882;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_0_5 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_0_5 <= _GEN_883;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_0_6 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_0_6 <= _GEN_884;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_0_7 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_0_7 <= _GEN_885;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_0_8 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_0_8 <= _GEN_886;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_0_9 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_0_9 <= _GEN_887;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_0_10 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_0_10 <= _GEN_888;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_0_11 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_0_11 <= _GEN_889;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_0_12 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_0_12 <= _GEN_890;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_0_13 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_0_13 <= _GEN_891;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_0_14 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_0_14 <= _GEN_892;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_0_15 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_0_15 <= _GEN_893;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_1_0 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_1_0 <= _GEN_894;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_1_1 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_1_1 <= _GEN_895;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_1_2 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_1_2 <= _GEN_896;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_1_3 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_1_3 <= _GEN_897;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_1_4 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_1_4 <= _GEN_898;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_1_5 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_1_5 <= _GEN_899;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_1_6 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_1_6 <= _GEN_900;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_1_7 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_1_7 <= _GEN_901;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_1_8 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_1_8 <= _GEN_902;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_1_9 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_1_9 <= _GEN_903;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_1_10 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_1_10 <= _GEN_904;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_1_11 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_1_11 <= _GEN_905;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_1_12 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_1_12 <= _GEN_906;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_1_13 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_1_13 <= _GEN_907;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_1_14 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_1_14 <= _GEN_908;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_1_15 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_1_15 <= _GEN_909;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_2_0 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_2_0 <= _GEN_910;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_2_1 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_2_1 <= _GEN_911;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_2_2 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_2_2 <= _GEN_912;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_2_3 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_2_3 <= _GEN_913;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_2_4 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_2_4 <= _GEN_914;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_2_5 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_2_5 <= _GEN_915;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_2_6 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_2_6 <= _GEN_916;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_2_7 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_2_7 <= _GEN_917;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_2_8 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_2_8 <= _GEN_918;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_2_9 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_2_9 <= _GEN_919;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_2_10 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_2_10 <= _GEN_920;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_2_11 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_2_11 <= _GEN_921;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_2_12 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_2_12 <= _GEN_922;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_2_13 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_2_13 <= _GEN_923;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_2_14 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_2_14 <= _GEN_924;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_2_15 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_2_15 <= _GEN_925;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_3_0 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_3_0 <= _GEN_926;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_3_1 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_3_1 <= _GEN_927;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_3_2 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_3_2 <= _GEN_928;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_3_3 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_3_3 <= _GEN_929;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_3_4 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_3_4 <= _GEN_930;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_3_5 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_3_5 <= _GEN_931;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_3_6 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_3_6 <= _GEN_932;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_3_7 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_3_7 <= _GEN_933;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_3_8 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_3_8 <= _GEN_934;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_3_9 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_3_9 <= _GEN_935;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_3_10 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_3_10 <= _GEN_936;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_3_11 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_3_11 <= _GEN_937;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_3_12 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_3_12 <= _GEN_938;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_3_13 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_3_13 <= _GEN_939;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_3_14 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_3_14 <= _GEN_940;
        end
      end
    end
    if (reset) begin // @[dcache.scala 92:26]
      tag_3_15 <= 22'h0; // @[dcache.scala 92:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          tag_3_15 <= _GEN_941;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_0_0 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_0_0 <= _GEN_942;
        end else begin
          valid_0_0 <= _GEN_1751;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_0_1 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_0_1 <= _GEN_943;
        end else begin
          valid_0_1 <= _GEN_1752;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_0_2 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_0_2 <= _GEN_944;
        end else begin
          valid_0_2 <= _GEN_1753;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_0_3 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_0_3 <= _GEN_945;
        end else begin
          valid_0_3 <= _GEN_1754;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_0_4 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_0_4 <= _GEN_946;
        end else begin
          valid_0_4 <= _GEN_1755;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_0_5 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_0_5 <= _GEN_947;
        end else begin
          valid_0_5 <= _GEN_1756;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_0_6 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_0_6 <= _GEN_948;
        end else begin
          valid_0_6 <= _GEN_1757;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_0_7 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_0_7 <= _GEN_949;
        end else begin
          valid_0_7 <= _GEN_1758;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_0_8 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_0_8 <= _GEN_950;
        end else begin
          valid_0_8 <= _GEN_1759;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_0_9 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_0_9 <= _GEN_951;
        end else begin
          valid_0_9 <= _GEN_1760;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_0_10 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_0_10 <= _GEN_952;
        end else begin
          valid_0_10 <= _GEN_1761;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_0_11 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_0_11 <= _GEN_953;
        end else begin
          valid_0_11 <= _GEN_1762;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_0_12 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_0_12 <= _GEN_954;
        end else begin
          valid_0_12 <= _GEN_1763;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_0_13 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_0_13 <= _GEN_955;
        end else begin
          valid_0_13 <= _GEN_1764;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_0_14 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_0_14 <= _GEN_956;
        end else begin
          valid_0_14 <= _GEN_1765;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_0_15 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_0_15 <= _GEN_957;
        end else begin
          valid_0_15 <= _GEN_1766;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_1_0 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_1_0 <= _GEN_958;
        end else begin
          valid_1_0 <= _GEN_1767;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_1_1 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_1_1 <= _GEN_959;
        end else begin
          valid_1_1 <= _GEN_1768;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_1_2 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_1_2 <= _GEN_960;
        end else begin
          valid_1_2 <= _GEN_1769;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_1_3 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_1_3 <= _GEN_961;
        end else begin
          valid_1_3 <= _GEN_1770;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_1_4 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_1_4 <= _GEN_962;
        end else begin
          valid_1_4 <= _GEN_1771;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_1_5 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_1_5 <= _GEN_963;
        end else begin
          valid_1_5 <= _GEN_1772;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_1_6 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_1_6 <= _GEN_964;
        end else begin
          valid_1_6 <= _GEN_1773;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_1_7 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_1_7 <= _GEN_965;
        end else begin
          valid_1_7 <= _GEN_1774;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_1_8 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_1_8 <= _GEN_966;
        end else begin
          valid_1_8 <= _GEN_1775;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_1_9 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_1_9 <= _GEN_967;
        end else begin
          valid_1_9 <= _GEN_1776;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_1_10 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_1_10 <= _GEN_968;
        end else begin
          valid_1_10 <= _GEN_1777;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_1_11 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_1_11 <= _GEN_969;
        end else begin
          valid_1_11 <= _GEN_1778;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_1_12 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_1_12 <= _GEN_970;
        end else begin
          valid_1_12 <= _GEN_1779;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_1_13 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_1_13 <= _GEN_971;
        end else begin
          valid_1_13 <= _GEN_1780;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_1_14 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_1_14 <= _GEN_972;
        end else begin
          valid_1_14 <= _GEN_1781;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_1_15 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_1_15 <= _GEN_973;
        end else begin
          valid_1_15 <= _GEN_1782;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_2_0 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_2_0 <= _GEN_974;
        end else begin
          valid_2_0 <= _GEN_1783;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_2_1 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_2_1 <= _GEN_975;
        end else begin
          valid_2_1 <= _GEN_1784;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_2_2 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_2_2 <= _GEN_976;
        end else begin
          valid_2_2 <= _GEN_1785;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_2_3 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_2_3 <= _GEN_977;
        end else begin
          valid_2_3 <= _GEN_1786;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_2_4 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_2_4 <= _GEN_978;
        end else begin
          valid_2_4 <= _GEN_1787;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_2_5 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_2_5 <= _GEN_979;
        end else begin
          valid_2_5 <= _GEN_1788;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_2_6 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_2_6 <= _GEN_980;
        end else begin
          valid_2_6 <= _GEN_1789;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_2_7 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_2_7 <= _GEN_981;
        end else begin
          valid_2_7 <= _GEN_1790;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_2_8 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_2_8 <= _GEN_982;
        end else begin
          valid_2_8 <= _GEN_1791;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_2_9 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_2_9 <= _GEN_983;
        end else begin
          valid_2_9 <= _GEN_1792;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_2_10 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_2_10 <= _GEN_984;
        end else begin
          valid_2_10 <= _GEN_1793;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_2_11 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_2_11 <= _GEN_985;
        end else begin
          valid_2_11 <= _GEN_1794;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_2_12 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_2_12 <= _GEN_986;
        end else begin
          valid_2_12 <= _GEN_1795;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_2_13 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_2_13 <= _GEN_987;
        end else begin
          valid_2_13 <= _GEN_1796;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_2_14 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_2_14 <= _GEN_988;
        end else begin
          valid_2_14 <= _GEN_1797;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_2_15 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_2_15 <= _GEN_989;
        end else begin
          valid_2_15 <= _GEN_1798;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_3_0 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_3_0 <= _GEN_990;
        end else begin
          valid_3_0 <= _GEN_1799;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_3_1 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_3_1 <= _GEN_991;
        end else begin
          valid_3_1 <= _GEN_1800;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_3_2 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_3_2 <= _GEN_992;
        end else begin
          valid_3_2 <= _GEN_1801;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_3_3 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_3_3 <= _GEN_993;
        end else begin
          valid_3_3 <= _GEN_1802;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_3_4 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_3_4 <= _GEN_994;
        end else begin
          valid_3_4 <= _GEN_1803;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_3_5 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_3_5 <= _GEN_995;
        end else begin
          valid_3_5 <= _GEN_1804;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_3_6 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_3_6 <= _GEN_996;
        end else begin
          valid_3_6 <= _GEN_1805;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_3_7 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_3_7 <= _GEN_997;
        end else begin
          valid_3_7 <= _GEN_1806;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_3_8 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_3_8 <= _GEN_998;
        end else begin
          valid_3_8 <= _GEN_1807;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_3_9 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_3_9 <= _GEN_999;
        end else begin
          valid_3_9 <= _GEN_1808;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_3_10 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_3_10 <= _GEN_1000;
        end else begin
          valid_3_10 <= _GEN_1809;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_3_11 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_3_11 <= _GEN_1001;
        end else begin
          valid_3_11 <= _GEN_1810;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_3_12 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_3_12 <= _GEN_1002;
        end else begin
          valid_3_12 <= _GEN_1811;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_3_13 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_3_13 <= _GEN_1003;
        end else begin
          valid_3_13 <= _GEN_1812;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_3_14 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_3_14 <= _GEN_1004;
        end else begin
          valid_3_14 <= _GEN_1813;
        end
      end
    end
    if (reset) begin // @[dcache.scala 93:26]
      valid_3_15 <= 1'h0; // @[dcache.scala 93:26]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          valid_3_15 <= _GEN_1005;
        end else begin
          valid_3_15 <= _GEN_1814;
        end
      end
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_0_0 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_0_0 <= _GEN_390;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_0_0 <= _GEN_390;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_0_0 <= _GEN_390;
    end else begin
      dirty_0_0 <= _GEN_1815;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_0_1 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_0_1 <= _GEN_391;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_0_1 <= _GEN_391;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_0_1 <= _GEN_391;
    end else begin
      dirty_0_1 <= _GEN_1816;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_0_2 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_0_2 <= _GEN_392;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_0_2 <= _GEN_392;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_0_2 <= _GEN_392;
    end else begin
      dirty_0_2 <= _GEN_1817;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_0_3 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_0_3 <= _GEN_393;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_0_3 <= _GEN_393;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_0_3 <= _GEN_393;
    end else begin
      dirty_0_3 <= _GEN_1818;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_0_4 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_0_4 <= _GEN_394;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_0_4 <= _GEN_394;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_0_4 <= _GEN_394;
    end else begin
      dirty_0_4 <= _GEN_1819;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_0_5 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_0_5 <= _GEN_395;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_0_5 <= _GEN_395;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_0_5 <= _GEN_395;
    end else begin
      dirty_0_5 <= _GEN_1820;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_0_6 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_0_6 <= _GEN_396;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_0_6 <= _GEN_396;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_0_6 <= _GEN_396;
    end else begin
      dirty_0_6 <= _GEN_1821;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_0_7 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_0_7 <= _GEN_397;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_0_7 <= _GEN_397;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_0_7 <= _GEN_397;
    end else begin
      dirty_0_7 <= _GEN_1822;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_0_8 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_0_8 <= _GEN_398;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_0_8 <= _GEN_398;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_0_8 <= _GEN_398;
    end else begin
      dirty_0_8 <= _GEN_1823;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_0_9 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_0_9 <= _GEN_399;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_0_9 <= _GEN_399;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_0_9 <= _GEN_399;
    end else begin
      dirty_0_9 <= _GEN_1824;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_0_10 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_0_10 <= _GEN_400;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_0_10 <= _GEN_400;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_0_10 <= _GEN_400;
    end else begin
      dirty_0_10 <= _GEN_1825;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_0_11 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_0_11 <= _GEN_401;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_0_11 <= _GEN_401;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_0_11 <= _GEN_401;
    end else begin
      dirty_0_11 <= _GEN_1826;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_0_12 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_0_12 <= _GEN_402;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_0_12 <= _GEN_402;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_0_12 <= _GEN_402;
    end else begin
      dirty_0_12 <= _GEN_1827;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_0_13 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_0_13 <= _GEN_403;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_0_13 <= _GEN_403;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_0_13 <= _GEN_403;
    end else begin
      dirty_0_13 <= _GEN_1828;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_0_14 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_0_14 <= _GEN_404;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_0_14 <= _GEN_404;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_0_14 <= _GEN_404;
    end else begin
      dirty_0_14 <= _GEN_1829;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_0_15 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_0_15 <= _GEN_405;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_0_15 <= _GEN_405;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_0_15 <= _GEN_405;
    end else begin
      dirty_0_15 <= _GEN_1830;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_1_0 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_1_0 <= _GEN_406;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_1_0 <= _GEN_406;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_1_0 <= _GEN_406;
    end else begin
      dirty_1_0 <= _GEN_1831;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_1_1 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_1_1 <= _GEN_407;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_1_1 <= _GEN_407;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_1_1 <= _GEN_407;
    end else begin
      dirty_1_1 <= _GEN_1832;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_1_2 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_1_2 <= _GEN_408;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_1_2 <= _GEN_408;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_1_2 <= _GEN_408;
    end else begin
      dirty_1_2 <= _GEN_1833;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_1_3 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_1_3 <= _GEN_409;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_1_3 <= _GEN_409;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_1_3 <= _GEN_409;
    end else begin
      dirty_1_3 <= _GEN_1834;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_1_4 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_1_4 <= _GEN_410;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_1_4 <= _GEN_410;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_1_4 <= _GEN_410;
    end else begin
      dirty_1_4 <= _GEN_1835;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_1_5 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_1_5 <= _GEN_411;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_1_5 <= _GEN_411;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_1_5 <= _GEN_411;
    end else begin
      dirty_1_5 <= _GEN_1836;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_1_6 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_1_6 <= _GEN_412;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_1_6 <= _GEN_412;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_1_6 <= _GEN_412;
    end else begin
      dirty_1_6 <= _GEN_1837;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_1_7 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_1_7 <= _GEN_413;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_1_7 <= _GEN_413;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_1_7 <= _GEN_413;
    end else begin
      dirty_1_7 <= _GEN_1838;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_1_8 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_1_8 <= _GEN_414;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_1_8 <= _GEN_414;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_1_8 <= _GEN_414;
    end else begin
      dirty_1_8 <= _GEN_1839;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_1_9 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_1_9 <= _GEN_415;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_1_9 <= _GEN_415;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_1_9 <= _GEN_415;
    end else begin
      dirty_1_9 <= _GEN_1840;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_1_10 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_1_10 <= _GEN_416;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_1_10 <= _GEN_416;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_1_10 <= _GEN_416;
    end else begin
      dirty_1_10 <= _GEN_1841;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_1_11 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_1_11 <= _GEN_417;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_1_11 <= _GEN_417;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_1_11 <= _GEN_417;
    end else begin
      dirty_1_11 <= _GEN_1842;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_1_12 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_1_12 <= _GEN_418;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_1_12 <= _GEN_418;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_1_12 <= _GEN_418;
    end else begin
      dirty_1_12 <= _GEN_1843;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_1_13 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_1_13 <= _GEN_419;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_1_13 <= _GEN_419;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_1_13 <= _GEN_419;
    end else begin
      dirty_1_13 <= _GEN_1844;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_1_14 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_1_14 <= _GEN_420;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_1_14 <= _GEN_420;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_1_14 <= _GEN_420;
    end else begin
      dirty_1_14 <= _GEN_1845;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_1_15 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_1_15 <= _GEN_421;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_1_15 <= _GEN_421;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_1_15 <= _GEN_421;
    end else begin
      dirty_1_15 <= _GEN_1846;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_2_0 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_2_0 <= _GEN_422;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_2_0 <= _GEN_422;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_2_0 <= _GEN_422;
    end else begin
      dirty_2_0 <= _GEN_1847;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_2_1 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_2_1 <= _GEN_423;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_2_1 <= _GEN_423;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_2_1 <= _GEN_423;
    end else begin
      dirty_2_1 <= _GEN_1848;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_2_2 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_2_2 <= _GEN_424;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_2_2 <= _GEN_424;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_2_2 <= _GEN_424;
    end else begin
      dirty_2_2 <= _GEN_1849;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_2_3 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_2_3 <= _GEN_425;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_2_3 <= _GEN_425;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_2_3 <= _GEN_425;
    end else begin
      dirty_2_3 <= _GEN_1850;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_2_4 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_2_4 <= _GEN_426;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_2_4 <= _GEN_426;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_2_4 <= _GEN_426;
    end else begin
      dirty_2_4 <= _GEN_1851;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_2_5 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_2_5 <= _GEN_427;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_2_5 <= _GEN_427;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_2_5 <= _GEN_427;
    end else begin
      dirty_2_5 <= _GEN_1852;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_2_6 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_2_6 <= _GEN_428;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_2_6 <= _GEN_428;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_2_6 <= _GEN_428;
    end else begin
      dirty_2_6 <= _GEN_1853;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_2_7 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_2_7 <= _GEN_429;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_2_7 <= _GEN_429;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_2_7 <= _GEN_429;
    end else begin
      dirty_2_7 <= _GEN_1854;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_2_8 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_2_8 <= _GEN_430;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_2_8 <= _GEN_430;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_2_8 <= _GEN_430;
    end else begin
      dirty_2_8 <= _GEN_1855;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_2_9 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_2_9 <= _GEN_431;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_2_9 <= _GEN_431;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_2_9 <= _GEN_431;
    end else begin
      dirty_2_9 <= _GEN_1856;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_2_10 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_2_10 <= _GEN_432;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_2_10 <= _GEN_432;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_2_10 <= _GEN_432;
    end else begin
      dirty_2_10 <= _GEN_1857;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_2_11 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_2_11 <= _GEN_433;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_2_11 <= _GEN_433;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_2_11 <= _GEN_433;
    end else begin
      dirty_2_11 <= _GEN_1858;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_2_12 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_2_12 <= _GEN_434;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_2_12 <= _GEN_434;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_2_12 <= _GEN_434;
    end else begin
      dirty_2_12 <= _GEN_1859;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_2_13 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_2_13 <= _GEN_435;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_2_13 <= _GEN_435;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_2_13 <= _GEN_435;
    end else begin
      dirty_2_13 <= _GEN_1860;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_2_14 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_2_14 <= _GEN_436;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_2_14 <= _GEN_436;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_2_14 <= _GEN_436;
    end else begin
      dirty_2_14 <= _GEN_1861;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_2_15 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_2_15 <= _GEN_437;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_2_15 <= _GEN_437;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_2_15 <= _GEN_437;
    end else begin
      dirty_2_15 <= _GEN_1862;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_3_0 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_3_0 <= _GEN_438;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_3_0 <= _GEN_438;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_3_0 <= _GEN_438;
    end else begin
      dirty_3_0 <= _GEN_1863;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_3_1 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_3_1 <= _GEN_439;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_3_1 <= _GEN_439;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_3_1 <= _GEN_439;
    end else begin
      dirty_3_1 <= _GEN_1864;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_3_2 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_3_2 <= _GEN_440;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_3_2 <= _GEN_440;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_3_2 <= _GEN_440;
    end else begin
      dirty_3_2 <= _GEN_1865;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_3_3 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_3_3 <= _GEN_441;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_3_3 <= _GEN_441;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_3_3 <= _GEN_441;
    end else begin
      dirty_3_3 <= _GEN_1866;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_3_4 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_3_4 <= _GEN_442;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_3_4 <= _GEN_442;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_3_4 <= _GEN_442;
    end else begin
      dirty_3_4 <= _GEN_1867;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_3_5 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_3_5 <= _GEN_443;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_3_5 <= _GEN_443;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_3_5 <= _GEN_443;
    end else begin
      dirty_3_5 <= _GEN_1868;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_3_6 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_3_6 <= _GEN_444;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_3_6 <= _GEN_444;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_3_6 <= _GEN_444;
    end else begin
      dirty_3_6 <= _GEN_1869;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_3_7 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_3_7 <= _GEN_445;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_3_7 <= _GEN_445;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_3_7 <= _GEN_445;
    end else begin
      dirty_3_7 <= _GEN_1870;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_3_8 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_3_8 <= _GEN_446;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_3_8 <= _GEN_446;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_3_8 <= _GEN_446;
    end else begin
      dirty_3_8 <= _GEN_1871;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_3_9 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_3_9 <= _GEN_447;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_3_9 <= _GEN_447;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_3_9 <= _GEN_447;
    end else begin
      dirty_3_9 <= _GEN_1872;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_3_10 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_3_10 <= _GEN_448;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_3_10 <= _GEN_448;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_3_10 <= _GEN_448;
    end else begin
      dirty_3_10 <= _GEN_1873;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_3_11 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_3_11 <= _GEN_449;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_3_11 <= _GEN_449;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_3_11 <= _GEN_449;
    end else begin
      dirty_3_11 <= _GEN_1874;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_3_12 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_3_12 <= _GEN_450;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_3_12 <= _GEN_450;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_3_12 <= _GEN_450;
    end else begin
      dirty_3_12 <= _GEN_1875;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_3_13 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_3_13 <= _GEN_451;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_3_13 <= _GEN_451;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_3_13 <= _GEN_451;
    end else begin
      dirty_3_13 <= _GEN_1876;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_3_14 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_3_14 <= _GEN_452;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_3_14 <= _GEN_452;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_3_14 <= _GEN_452;
    end else begin
      dirty_3_14 <= _GEN_1877;
    end
    if (reset) begin // @[dcache.scala 94:26]
      dirty_3_15 <= 1'h0; // @[dcache.scala 94:26]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      dirty_3_15 <= _GEN_453;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      dirty_3_15 <= _GEN_453;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      dirty_3_15 <= _GEN_453;
    end else begin
      dirty_3_15 <= _GEN_1878;
    end
    if (reset) begin // @[dcache.scala 96:30]
      wait_r <= 1'h0; // @[dcache.scala 96:30]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      if (!(flush_r | io_flush)) begin // @[dcache.scala 229:38]
        if (!(~hs_in & _io_dcRW_ready_T)) begin // @[dcache.scala 231:42]
          wait_r <= _GEN_592;
        end
      end
    end else if (!(_T_74)) begin // @[Conditional.scala 39:67]
      if (!(_T_76)) begin // @[Conditional.scala 39:67]
        wait_r <= _GEN_1881;
      end
    end
    if (reset) begin // @[dcache.scala 97:30]
      valid_r <= 1'h0; // @[dcache.scala 97:30]
    end else begin
      valid_r <= _GEN_2295;
    end
    if (reset) begin // @[dcache.scala 98:30]
      flush_r <= 1'h0; // @[dcache.scala 98:30]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      flush_r <= _GEN_134;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      flush_r <= _GEN_134;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      flush_r <= _GEN_134;
    end else begin
      flush_r <= _GEN_1882;
    end
    if (reset) begin // @[dcache.scala 99:30]
      mode_r <= 5'h0; // @[dcache.scala 99:30]
    end else if (hs_in) begin // @[dcache.scala 120:16]
      mode_r <= io_dcRW_dc_mode; // @[dcache.scala 123:17]
    end
    if (reset) begin // @[dcache.scala 100:30]
      wdata_r <= 64'h0; // @[dcache.scala 100:30]
    end else if (hs_in) begin // @[dcache.scala 120:16]
      wdata_r <= io_dcRW_wdata; // @[dcache.scala 124:17]
    end
    if (reset) begin // @[dcache.scala 101:30]
      amo_r <= 5'h0; // @[dcache.scala 101:30]
    end else if (hs_in) begin // @[dcache.scala 120:16]
      amo_r <= io_dcRW_amo; // @[dcache.scala 125:17]
    end
    if (reset) begin // @[dcache.scala 108:34]
      addr_r <= 32'h0; // @[dcache.scala 108:34]
    end else if (hs_in) begin // @[dcache.scala 109:30]
      addr_r <= io_dcRW_addr;
    end
    if (reset) begin // @[dcache.scala 110:34]
      matchWay_r <= 2'h0; // @[dcache.scala 110:34]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      matchWay_r <= _GEN_129;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      matchWay_r <= _GEN_129;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      matchWay_r <= _GEN_129;
    end else begin
      matchWay_r <= _GEN_1883;
    end
    if (reset) begin // @[dcache.scala 111:34]
      offset <= 3'h0; // @[dcache.scala 111:34]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (_T_74) begin // @[Conditional.scala 39:67]
        offset <= 3'h0; // @[dcache.scala 257:20]
      end else if (_T_76) begin // @[Conditional.scala 39:67]
        offset <= _GEN_874;
      end else begin
        offset <= _GEN_1747;
      end
    end
    if (reset) begin // @[dcache.scala 112:34]
      rdatabuf <= 64'h0; // @[dcache.scala 112:34]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_76) begin // @[Conditional.scala 39:67]
          rdatabuf <= _GEN_876;
        end
      end
    end
    if (reset) begin // @[dcache.scala 114:34]
      blockIdx_r <= 4'h0; // @[dcache.scala 114:34]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      blockIdx_r <= _GEN_133;
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      blockIdx_r <= _GEN_133;
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      blockIdx_r <= _GEN_133;
    end else begin
      blockIdx_r <= _GEN_1884;
    end
    if (reset) begin // @[dcache.scala 153:24]
      state <= 3'h0; // @[dcache.scala 153:24]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      if (flush_r | io_flush) begin // @[dcache.scala 229:38]
        state <= 3'h6; // @[dcache.scala 230:23]
      end else if (!(~hs_in & _io_dcRW_ready_T)) begin // @[dcache.scala 231:42]
        state <= _GEN_590;
      end
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      if (axiRaddrEn & io_dataAxi_ra_ready) begin // @[dcache.scala 258:52]
        state <= 3'h2; // @[dcache.scala 259:25]
      end
    end else if (_T_76) begin // @[Conditional.scala 39:67]
      state <= _GEN_1006;
    end else begin
      state <= _GEN_1748;
    end
    if (reset) begin // @[dcache.scala 220:34]
      axiRdataEn <= 1'h0; // @[dcache.scala 220:34]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (_T_74) begin // @[Conditional.scala 39:67]
        axiRdataEn <= _GEN_613;
      end else if (_T_76) begin // @[Conditional.scala 39:67]
        axiRdataEn <= _GEN_877;
      end
    end
    if (reset) begin // @[dcache.scala 218:34]
      axiRaddrEn <= 1'h0; // @[dcache.scala 218:34]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      if (!(flush_r | io_flush)) begin // @[dcache.scala 229:38]
        if (!(~hs_in & _io_dcRW_ready_T)) begin // @[dcache.scala 231:42]
          axiRaddrEn <= _GEN_596;
        end
      end
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      if (axiRaddrEn & io_dataAxi_ra_ready) begin // @[dcache.scala 258:52]
        axiRaddrEn <= 1'h0; // @[dcache.scala 260:28]
      end
    end
    if (reset) begin // @[dcache.scala 221:34]
      axiWaddrEn <= 1'h0; // @[dcache.scala 221:34]
    end else if (_T_68) begin // @[Conditional.scala 40:58]
      if (!(flush_r | io_flush)) begin // @[dcache.scala 229:38]
        if (!(~hs_in & _io_dcRW_ready_T)) begin // @[dcache.scala 231:42]
          axiWaddrEn <= _GEN_595;
        end
      end
    end else if (!(_T_74)) begin // @[Conditional.scala 39:67]
      if (!(_T_76)) begin // @[Conditional.scala 39:67]
        axiWaddrEn <= _GEN_1749;
      end
    end
    if (reset) begin // @[dcache.scala 224:34]
      axiWdataEn <= 1'h0; // @[dcache.scala 224:34]
    end else if (!(_T_68)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (!(_T_76)) begin // @[Conditional.scala 39:67]
          axiWdataEn <= _GEN_1750;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_0_0 = _RAND_0[21:0];
  _RAND_1 = {1{`RANDOM}};
  tag_0_1 = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  tag_0_2 = _RAND_2[21:0];
  _RAND_3 = {1{`RANDOM}};
  tag_0_3 = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  tag_0_4 = _RAND_4[21:0];
  _RAND_5 = {1{`RANDOM}};
  tag_0_5 = _RAND_5[21:0];
  _RAND_6 = {1{`RANDOM}};
  tag_0_6 = _RAND_6[21:0];
  _RAND_7 = {1{`RANDOM}};
  tag_0_7 = _RAND_7[21:0];
  _RAND_8 = {1{`RANDOM}};
  tag_0_8 = _RAND_8[21:0];
  _RAND_9 = {1{`RANDOM}};
  tag_0_9 = _RAND_9[21:0];
  _RAND_10 = {1{`RANDOM}};
  tag_0_10 = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  tag_0_11 = _RAND_11[21:0];
  _RAND_12 = {1{`RANDOM}};
  tag_0_12 = _RAND_12[21:0];
  _RAND_13 = {1{`RANDOM}};
  tag_0_13 = _RAND_13[21:0];
  _RAND_14 = {1{`RANDOM}};
  tag_0_14 = _RAND_14[21:0];
  _RAND_15 = {1{`RANDOM}};
  tag_0_15 = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  tag_1_0 = _RAND_16[21:0];
  _RAND_17 = {1{`RANDOM}};
  tag_1_1 = _RAND_17[21:0];
  _RAND_18 = {1{`RANDOM}};
  tag_1_2 = _RAND_18[21:0];
  _RAND_19 = {1{`RANDOM}};
  tag_1_3 = _RAND_19[21:0];
  _RAND_20 = {1{`RANDOM}};
  tag_1_4 = _RAND_20[21:0];
  _RAND_21 = {1{`RANDOM}};
  tag_1_5 = _RAND_21[21:0];
  _RAND_22 = {1{`RANDOM}};
  tag_1_6 = _RAND_22[21:0];
  _RAND_23 = {1{`RANDOM}};
  tag_1_7 = _RAND_23[21:0];
  _RAND_24 = {1{`RANDOM}};
  tag_1_8 = _RAND_24[21:0];
  _RAND_25 = {1{`RANDOM}};
  tag_1_9 = _RAND_25[21:0];
  _RAND_26 = {1{`RANDOM}};
  tag_1_10 = _RAND_26[21:0];
  _RAND_27 = {1{`RANDOM}};
  tag_1_11 = _RAND_27[21:0];
  _RAND_28 = {1{`RANDOM}};
  tag_1_12 = _RAND_28[21:0];
  _RAND_29 = {1{`RANDOM}};
  tag_1_13 = _RAND_29[21:0];
  _RAND_30 = {1{`RANDOM}};
  tag_1_14 = _RAND_30[21:0];
  _RAND_31 = {1{`RANDOM}};
  tag_1_15 = _RAND_31[21:0];
  _RAND_32 = {1{`RANDOM}};
  tag_2_0 = _RAND_32[21:0];
  _RAND_33 = {1{`RANDOM}};
  tag_2_1 = _RAND_33[21:0];
  _RAND_34 = {1{`RANDOM}};
  tag_2_2 = _RAND_34[21:0];
  _RAND_35 = {1{`RANDOM}};
  tag_2_3 = _RAND_35[21:0];
  _RAND_36 = {1{`RANDOM}};
  tag_2_4 = _RAND_36[21:0];
  _RAND_37 = {1{`RANDOM}};
  tag_2_5 = _RAND_37[21:0];
  _RAND_38 = {1{`RANDOM}};
  tag_2_6 = _RAND_38[21:0];
  _RAND_39 = {1{`RANDOM}};
  tag_2_7 = _RAND_39[21:0];
  _RAND_40 = {1{`RANDOM}};
  tag_2_8 = _RAND_40[21:0];
  _RAND_41 = {1{`RANDOM}};
  tag_2_9 = _RAND_41[21:0];
  _RAND_42 = {1{`RANDOM}};
  tag_2_10 = _RAND_42[21:0];
  _RAND_43 = {1{`RANDOM}};
  tag_2_11 = _RAND_43[21:0];
  _RAND_44 = {1{`RANDOM}};
  tag_2_12 = _RAND_44[21:0];
  _RAND_45 = {1{`RANDOM}};
  tag_2_13 = _RAND_45[21:0];
  _RAND_46 = {1{`RANDOM}};
  tag_2_14 = _RAND_46[21:0];
  _RAND_47 = {1{`RANDOM}};
  tag_2_15 = _RAND_47[21:0];
  _RAND_48 = {1{`RANDOM}};
  tag_3_0 = _RAND_48[21:0];
  _RAND_49 = {1{`RANDOM}};
  tag_3_1 = _RAND_49[21:0];
  _RAND_50 = {1{`RANDOM}};
  tag_3_2 = _RAND_50[21:0];
  _RAND_51 = {1{`RANDOM}};
  tag_3_3 = _RAND_51[21:0];
  _RAND_52 = {1{`RANDOM}};
  tag_3_4 = _RAND_52[21:0];
  _RAND_53 = {1{`RANDOM}};
  tag_3_5 = _RAND_53[21:0];
  _RAND_54 = {1{`RANDOM}};
  tag_3_6 = _RAND_54[21:0];
  _RAND_55 = {1{`RANDOM}};
  tag_3_7 = _RAND_55[21:0];
  _RAND_56 = {1{`RANDOM}};
  tag_3_8 = _RAND_56[21:0];
  _RAND_57 = {1{`RANDOM}};
  tag_3_9 = _RAND_57[21:0];
  _RAND_58 = {1{`RANDOM}};
  tag_3_10 = _RAND_58[21:0];
  _RAND_59 = {1{`RANDOM}};
  tag_3_11 = _RAND_59[21:0];
  _RAND_60 = {1{`RANDOM}};
  tag_3_12 = _RAND_60[21:0];
  _RAND_61 = {1{`RANDOM}};
  tag_3_13 = _RAND_61[21:0];
  _RAND_62 = {1{`RANDOM}};
  tag_3_14 = _RAND_62[21:0];
  _RAND_63 = {1{`RANDOM}};
  tag_3_15 = _RAND_63[21:0];
  _RAND_64 = {1{`RANDOM}};
  valid_0_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_0_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_0_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  valid_0_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  valid_0_4 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  valid_0_5 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  valid_0_6 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  valid_0_7 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  valid_0_8 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  valid_0_9 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  valid_0_10 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid_0_11 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  valid_0_12 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  valid_0_13 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  valid_0_14 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  valid_0_15 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  valid_1_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_1_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_1_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_1_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_1_4 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_1_5 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_1_6 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_1_7 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_1_8 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_1_9 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_1_10 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_1_11 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_1_12 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_1_13 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_1_14 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_1_15 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  valid_2_0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  valid_2_1 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  valid_2_2 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  valid_2_3 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  valid_2_4 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  valid_2_5 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  valid_2_6 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  valid_2_7 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  valid_2_8 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  valid_2_9 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  valid_2_10 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  valid_2_11 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  valid_2_12 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  valid_2_13 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  valid_2_14 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  valid_2_15 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  valid_3_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  valid_3_1 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  valid_3_2 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  valid_3_3 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  valid_3_4 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  valid_3_5 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  valid_3_6 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  valid_3_7 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  valid_3_8 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  valid_3_9 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  valid_3_10 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  valid_3_11 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  valid_3_12 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  valid_3_13 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  valid_3_14 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  valid_3_15 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  dirty_0_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  dirty_0_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  dirty_0_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  dirty_0_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  dirty_0_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  dirty_0_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  dirty_0_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  dirty_0_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  dirty_0_8 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  dirty_0_9 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  dirty_0_10 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  dirty_0_11 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  dirty_0_12 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  dirty_0_13 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  dirty_0_14 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  dirty_0_15 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  dirty_1_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  dirty_1_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  dirty_1_2 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  dirty_1_3 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  dirty_1_4 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  dirty_1_5 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  dirty_1_6 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  dirty_1_7 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  dirty_1_8 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  dirty_1_9 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  dirty_1_10 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  dirty_1_11 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  dirty_1_12 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  dirty_1_13 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  dirty_1_14 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  dirty_1_15 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  dirty_2_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  dirty_2_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  dirty_2_2 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  dirty_2_3 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  dirty_2_4 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  dirty_2_5 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  dirty_2_6 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  dirty_2_7 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  dirty_2_8 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  dirty_2_9 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  dirty_2_10 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  dirty_2_11 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  dirty_2_12 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  dirty_2_13 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  dirty_2_14 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  dirty_2_15 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  dirty_3_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  dirty_3_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  dirty_3_2 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  dirty_3_3 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  dirty_3_4 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  dirty_3_5 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  dirty_3_6 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  dirty_3_7 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  dirty_3_8 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  dirty_3_9 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  dirty_3_10 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  dirty_3_11 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  dirty_3_12 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  dirty_3_13 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  dirty_3_14 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  dirty_3_15 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  wait_r = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  valid_r = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  flush_r = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  mode_r = _RAND_195[4:0];
  _RAND_196 = {2{`RANDOM}};
  wdata_r = _RAND_196[63:0];
  _RAND_197 = {1{`RANDOM}};
  amo_r = _RAND_197[4:0];
  _RAND_198 = {1{`RANDOM}};
  addr_r = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  matchWay_r = _RAND_199[1:0];
  _RAND_200 = {1{`RANDOM}};
  offset = _RAND_200[2:0];
  _RAND_201 = {2{`RANDOM}};
  rdatabuf = _RAND_201[63:0];
  _RAND_202 = {1{`RANDOM}};
  blockIdx_r = _RAND_202[3:0];
  _RAND_203 = {1{`RANDOM}};
  state = _RAND_203[2:0];
  _RAND_204 = {1{`RANDOM}};
  axiRdataEn = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  axiRaddrEn = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  axiWaddrEn = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  axiWdataEn = _RAND_207[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_ToAXI(
  input         clock,
  input         reset,
  input  [31:0] io_dataIO_addr,
  output [63:0] io_dataIO_rdata,
  output        io_dataIO_rvalid,
  input  [63:0] io_dataIO_wdata,
  input  [4:0]  io_dataIO_dc_mode,
  output        io_dataIO_ready,
  input         io_outAxi_wa_ready,
  output        io_outAxi_wa_valid,
  output [3:0]  io_outAxi_wa_bits_id,
  output [31:0] io_outAxi_wa_bits_addr,
  output [7:0]  io_outAxi_wa_bits_len,
  output [2:0]  io_outAxi_wa_bits_size,
  output [1:0]  io_outAxi_wa_bits_burst,
  input         io_outAxi_wd_ready,
  output        io_outAxi_wd_valid,
  output [63:0] io_outAxi_wd_bits_data,
  output [7:0]  io_outAxi_wd_bits_strb,
  output        io_outAxi_wd_bits_last,
  output        io_outAxi_wr_ready,
  input         io_outAxi_wr_valid,
  input  [3:0]  io_outAxi_wr_bits_id,
  input  [1:0]  io_outAxi_wr_bits_resp,
  input         io_outAxi_ra_ready,
  output        io_outAxi_ra_valid,
  output [3:0]  io_outAxi_ra_bits_id,
  output [31:0] io_outAxi_ra_bits_addr,
  output [7:0]  io_outAxi_ra_bits_len,
  output [2:0]  io_outAxi_ra_bits_size,
  output [1:0]  io_outAxi_ra_bits_burst,
  output        io_outAxi_rd_ready,
  input         io_outAxi_rd_valid,
  input  [3:0]  io_outAxi_rd_bits_id,
  input  [63:0] io_outAxi_rd_bits_data,
  input  [1:0]  io_outAxi_rd_bits_resp,
  input         io_outAxi_rd_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg  waddrEn; // @[toaxi.scala 66:26]
  reg [31:0] waddr; // @[toaxi.scala 67:26]
  reg [2:0] wsize; // @[toaxi.scala 68:26]
  reg  wdataEn; // @[toaxi.scala 71:26]
  reg [63:0] wdata; // @[toaxi.scala 72:26]
  reg [7:0] wstrb; // @[toaxi.scala 73:26]
  reg [2:0] rsize; // @[toaxi.scala 75:26]
  reg  raddrEn; // @[toaxi.scala 76:26]
  reg [31:0] raddr; // @[toaxi.scala 77:26]
  reg  rdataEn; // @[toaxi.scala 78:26]
  reg [63:0] rdata; // @[toaxi.scala 79:26]
  reg [31:0] pre_addr; // @[toaxi.scala 81:27]
  reg [4:0] mode; // @[toaxi.scala 85:23]
  reg [2:0] state; // @[toaxi.scala 92:25]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _wtype_T_1 = 5'h8 == io_dataIO_dc_mode; // @[Lookup.scala 31:38]
  wire  _wtype_T_3 = 5'h9 == io_dataIO_dc_mode; // @[Lookup.scala 31:38]
  wire  _wtype_T_5 = 5'ha == io_dataIO_dc_mode; // @[Lookup.scala 31:38]
  wire  _wtype_T_7 = 5'hb == io_dataIO_dc_mode; // @[Lookup.scala 31:38]
  wire [2:0] _wtype_T_8 = _wtype_T_7 ? 3'h3 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _wtype_T_9 = _wtype_T_5 ? 3'h2 : _wtype_T_8; // @[Lookup.scala 33:37]
  wire [2:0] _wtype_T_10 = _wtype_T_3 ? 3'h1 : _wtype_T_9; // @[Lookup.scala 33:37]
  wire [7:0] _wtype_T_11 = _wtype_T_7 ? 8'hff : 8'h0; // @[Lookup.scala 33:37]
  wire [7:0] _wtype_T_12 = _wtype_T_5 ? 8'hf : _wtype_T_11; // @[Lookup.scala 33:37]
  wire [7:0] _wtype_T_13 = _wtype_T_3 ? 8'h3 : _wtype_T_12; // @[Lookup.scala 33:37]
  wire [7:0] wtype_1 = _wtype_T_1 ? 8'h1 : _wtype_T_13; // @[Lookup.scala 33:37]
  wire [14:0] _GEN_84 = {{7'd0}, wtype_1}; // @[toaxi.scala 113:37]
  wire [14:0] _wstrb_T_1 = _GEN_84 << io_dataIO_addr[2:0]; // @[toaxi.scala 113:37]
  wire [6:0] _wdata_T_1 = io_dataIO_addr[2:0] * 4'h8; // @[toaxi.scala 114:55]
  wire [190:0] _GEN_85 = {{127'd0}, io_dataIO_wdata}; // @[toaxi.scala 114:38]
  wire [190:0] _wdata_T_2 = _GEN_85 << _wdata_T_1; // @[toaxi.scala 114:38]
  wire [2:0] _rsize_T_5 = 5'h5 == io_dataIO_dc_mode ? 3'h1 : 3'h0; // @[Mux.scala 80:57]
  wire [2:0] _rsize_T_7 = 5'h15 == io_dataIO_dc_mode ? 3'h1 : _rsize_T_5; // @[Mux.scala 80:57]
  wire [2:0] _rsize_T_9 = 5'h6 == io_dataIO_dc_mode ? 3'h2 : _rsize_T_7; // @[Mux.scala 80:57]
  wire [2:0] _rsize_T_11 = 5'h16 == io_dataIO_dc_mode ? 3'h2 : _rsize_T_9; // @[Mux.scala 80:57]
  wire [2:0] _rsize_T_13 = 5'h7 == io_dataIO_dc_mode ? 3'h3 : _rsize_T_11; // @[Mux.scala 80:57]
  wire  _GEN_4 = io_dataIO_dc_mode[2] | raddrEn; // @[toaxi.scala 116:43 toaxi.scala 130:25 toaxi.scala 76:26]
  wire  _GEN_8 = io_dataIO_dc_mode[3] | waddrEn; // @[toaxi.scala 101:37 toaxi.scala 105:25 toaxi.scala 66:26]
  wire [14:0] _GEN_10 = io_dataIO_dc_mode[3] ? _wstrb_T_1 : {{7'd0}, wstrb}; // @[toaxi.scala 101:37 toaxi.scala 113:25 toaxi.scala 73:26]
  wire  _T_6 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_8 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_21 = io_outAxi_wd_ready ? 3'h3 : state; // @[toaxi.scala 144:37 toaxi.scala 92:25]
  wire  _T_9 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_10 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _GEN_22 = raddrEn & io_outAxi_ra_ready ? 1'h0 : raddrEn; // @[toaxi.scala 157:48 toaxi.scala 158:25 toaxi.scala 76:26]
  wire [2:0] _GEN_24 = raddrEn & io_outAxi_ra_ready ? 3'h5 : state; // @[toaxi.scala 157:48 toaxi.scala 160:25 toaxi.scala 92:25]
  wire  _T_12 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire [2:0] strb_offset = pre_addr[2:0]; // @[toaxi.scala 169:43]
  wire  _T_14 = 5'h4 == mode; // @[Conditional.scala 37:30]
  wire [6:0] _tem_rdata_T = 4'h8 * strb_offset; // @[toaxi.scala 172:72]
  wire [63:0] _tem_rdata_T_1 = io_outAxi_rd_bits_data >> _tem_rdata_T; // @[toaxi.scala 172:64]
  wire [7:0] _tem_rdata_T_3 = _tem_rdata_T_1[7:0]; // @[toaxi.scala 172:94]
  wire  _T_15 = 5'h5 == mode; // @[Conditional.scala 37:30]
  wire [15:0] _tem_rdata_T_7 = _tem_rdata_T_1[15:0]; // @[toaxi.scala 176:95]
  wire  _T_16 = 5'h6 == mode; // @[Conditional.scala 37:30]
  wire [31:0] _tem_rdata_T_11 = _tem_rdata_T_1[31:0]; // @[toaxi.scala 180:95]
  wire [31:0] _GEN_29 = _T_16 ? $signed(_tem_rdata_T_11) : $signed(32'sh0); // @[Conditional.scala 39:67 toaxi.scala 180:37 toaxi.scala 168:29]
  wire [31:0] _GEN_31 = _T_15 ? $signed({{16{_tem_rdata_T_7[15]}},_tem_rdata_T_7}) : $signed(_GEN_29); // @[Conditional.scala 39:67 toaxi.scala 176:37]
  wire [31:0] _GEN_33 = _T_14 ? $signed({{24{_tem_rdata_T_3[7]}},_tem_rdata_T_3}) : $signed(_GEN_31); // @[Conditional.scala 40:58 toaxi.scala 172:37]
  wire [63:0] _rdata_T = {{32{_GEN_33[31]}},_GEN_33}; // @[toaxi.scala 173:50]
  wire  _T_17 = 5'h7 == mode; // @[Conditional.scala 37:30]
  wire  _T_18 = 5'h14 == mode; // @[Conditional.scala 37:30]
  wire  _T_19 = 5'h15 == mode; // @[Conditional.scala 37:30]
  wire  _T_20 = 5'h16 == mode; // @[Conditional.scala 37:30]
  wire [63:0] _GEN_25 = _T_20 ? {{32'd0}, _tem_rdata_T_1[31:0]} : rdata; // @[Conditional.scala 39:67 toaxi.scala 193:33 toaxi.scala 79:26]
  wire [63:0] _GEN_26 = _T_19 ? {{48'd0}, _tem_rdata_T_1[15:0]} : _GEN_25; // @[Conditional.scala 39:67 toaxi.scala 190:33]
  wire [63:0] _GEN_27 = _T_18 ? {{56'd0}, _tem_rdata_T_1[7:0]} : _GEN_26; // @[Conditional.scala 39:67 toaxi.scala 187:33]
  wire [63:0] _GEN_28 = _T_17 ? io_outAxi_rd_bits_data : _GEN_27; // @[Conditional.scala 39:67 toaxi.scala 184:37]
  wire [63:0] _GEN_30 = _T_16 ? _rdata_T : _GEN_28; // @[Conditional.scala 39:67 toaxi.scala 181:37]
  wire [63:0] _GEN_32 = _T_15 ? _rdata_T : _GEN_30; // @[Conditional.scala 39:67 toaxi.scala 177:37]
  wire [63:0] _GEN_34 = _T_14 ? _rdata_T : _GEN_32; // @[Conditional.scala 40:58 toaxi.scala 173:37]
  wire [63:0] _GEN_35 = rdataEn & io_outAxi_rd_valid ? _GEN_34 : rdata; // @[toaxi.scala 166:48 toaxi.scala 79:26]
  wire  _GEN_37 = rdataEn & io_outAxi_rd_valid ? 1'h0 : 1'h1; // @[toaxi.scala 166:48 toaxi.scala 198:25 toaxi.scala 164:21]
  wire [2:0] _GEN_38 = rdataEn & io_outAxi_rd_valid ? 3'h6 : state; // @[toaxi.scala 166:48 toaxi.scala 199:25 toaxi.scala 92:25]
  wire  _T_21 = 3'h6 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_39 = _T_21 ? 3'h0 : state; // @[Conditional.scala 39:67 toaxi.scala 203:19 toaxi.scala 92:25]
  wire  _GEN_40 = _T_12 ? _GEN_37 : rdataEn; // @[Conditional.scala 39:67 toaxi.scala 78:26]
  wire [63:0] _GEN_41 = _T_12 ? _GEN_35 : rdata; // @[Conditional.scala 39:67 toaxi.scala 79:26]
  wire [2:0] _GEN_43 = _T_12 ? _GEN_38 : _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_44 = _T_10 ? _GEN_22 : raddrEn; // @[Conditional.scala 39:67 toaxi.scala 76:26]
  wire [2:0] _GEN_46 = _T_10 ? _GEN_24 : _GEN_43; // @[Conditional.scala 39:67]
  wire  _GEN_47 = _T_10 ? rdataEn : _GEN_40; // @[Conditional.scala 39:67 toaxi.scala 78:26]
  wire [63:0] _GEN_48 = _T_10 ? rdata : _GEN_41; // @[Conditional.scala 39:67 toaxi.scala 79:26]
  wire  _GEN_49 = _T_9 ? 1'h0 : wdataEn; // @[Conditional.scala 39:67 toaxi.scala 152:21 toaxi.scala 71:26]
  wire [2:0] _GEN_50 = _T_9 ? 3'h0 : _GEN_46; // @[Conditional.scala 39:67 toaxi.scala 153:21]
  wire  _GEN_51 = _T_9 ? raddrEn : _GEN_44; // @[Conditional.scala 39:67 toaxi.scala 76:26]
  wire  _GEN_53 = _T_9 ? rdataEn : _GEN_47; // @[Conditional.scala 39:67 toaxi.scala 78:26]
  wire [63:0] _GEN_54 = _T_9 ? rdata : _GEN_48; // @[Conditional.scala 39:67 toaxi.scala 79:26]
  wire  _GEN_55 = _T_8 | _GEN_49; // @[Conditional.scala 39:67 toaxi.scala 143:21]
  wire [14:0] _GEN_74 = _T ? _GEN_10 : {{7'd0}, wstrb}; // @[Conditional.scala 40:58 toaxi.scala 73:26]
  reg [63:0] out_rdata; // @[toaxi.scala 208:28]
  reg  out_valid; // @[toaxi.scala 209:28]
  assign io_dataIO_rdata = out_rdata; // @[toaxi.scala 213:25]
  assign io_dataIO_rvalid = out_valid; // @[toaxi.scala 212:25]
  assign io_dataIO_ready = state == 3'h0; // @[toaxi.scala 206:31]
  assign io_outAxi_wa_valid = waddrEn; // @[toaxi.scala 217:31]
  assign io_outAxi_wa_bits_id = 4'h0; // @[axi.scala 41:38 axi.scala 41:38]
  assign io_outAxi_wa_bits_addr = waddr; // @[toaxi.scala 218:31]
  assign io_outAxi_wa_bits_len = 8'h0; // @[toaxi.scala 219:31]
  assign io_outAxi_wa_bits_size = wsize; // @[toaxi.scala 220:31]
  assign io_outAxi_wa_bits_burst = 2'h1; // @[toaxi.scala 221:31]
  assign io_outAxi_wd_valid = wdataEn; // @[toaxi.scala 223:31]
  assign io_outAxi_wd_bits_data = wdata; // @[toaxi.scala 224:31]
  assign io_outAxi_wd_bits_strb = wstrb; // @[toaxi.scala 225:31]
  assign io_outAxi_wd_bits_last = 1'h1; // @[toaxi.scala 70:27]
  assign io_outAxi_wr_ready = 1'h1; // @[toaxi.scala 228:31]
  assign io_outAxi_ra_valid = raddrEn; // @[toaxi.scala 230:31]
  assign io_outAxi_ra_bits_id = 4'h0; // @[axi.scala 41:38 axi.scala 41:38]
  assign io_outAxi_ra_bits_addr = raddr; // @[toaxi.scala 231:31]
  assign io_outAxi_ra_bits_len = 8'h0; // @[toaxi.scala 232:31]
  assign io_outAxi_ra_bits_size = rsize; // @[toaxi.scala 233:31]
  assign io_outAxi_ra_bits_burst = 2'h1; // @[toaxi.scala 234:31]
  assign io_outAxi_rd_ready = rdataEn; // @[toaxi.scala 236:31]
  always @(posedge clock) begin
    if (reset) begin // @[toaxi.scala 66:26]
      waddrEn <= 1'h0; // @[toaxi.scala 66:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      waddrEn <= _GEN_8;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      if (waddrEn & io_outAxi_wa_ready) begin // @[toaxi.scala 136:48]
        waddrEn <= 1'h0; // @[toaxi.scala 137:25]
      end
    end
    if (reset) begin // @[toaxi.scala 67:26]
      waddr <= 32'h0; // @[toaxi.scala 67:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_dataIO_dc_mode[3]) begin // @[toaxi.scala 101:37]
        waddr <= io_dataIO_addr; // @[toaxi.scala 103:25]
      end
    end
    if (reset) begin // @[toaxi.scala 68:26]
      wsize <= 3'h0; // @[toaxi.scala 68:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_dataIO_dc_mode[3]) begin // @[toaxi.scala 101:37]
        if (_wtype_T_1) begin // @[Lookup.scala 33:37]
          wsize <= 3'h0;
        end else begin
          wsize <= _wtype_T_10;
        end
      end
    end
    if (reset) begin // @[toaxi.scala 71:26]
      wdataEn <= 1'h0; // @[toaxi.scala 71:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_6)) begin // @[Conditional.scala 39:67]
        wdataEn <= _GEN_55;
      end
    end
    if (reset) begin // @[toaxi.scala 72:26]
      wdata <= 64'h0; // @[toaxi.scala 72:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_dataIO_dc_mode[3]) begin // @[toaxi.scala 101:37]
        wdata <= _wdata_T_2[63:0]; // @[toaxi.scala 114:25]
      end
    end
    if (reset) begin // @[toaxi.scala 73:26]
      wstrb <= 8'h0; // @[toaxi.scala 73:26]
    end else begin
      wstrb <= _GEN_74[7:0];
    end
    if (reset) begin // @[toaxi.scala 75:26]
      rsize <= 3'h0; // @[toaxi.scala 75:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (!(io_dataIO_dc_mode[3])) begin // @[toaxi.scala 101:37]
        if (io_dataIO_dc_mode[2]) begin // @[toaxi.scala 116:43]
          rsize <= _rsize_T_13; // @[toaxi.scala 118:23]
        end
      end
    end
    if (reset) begin // @[toaxi.scala 76:26]
      raddrEn <= 1'h0; // @[toaxi.scala 76:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (!(io_dataIO_dc_mode[3])) begin // @[toaxi.scala 101:37]
        raddrEn <= _GEN_4;
      end
    end else if (!(_T_6)) begin // @[Conditional.scala 39:67]
      if (!(_T_8)) begin // @[Conditional.scala 39:67]
        raddrEn <= _GEN_51;
      end
    end
    if (reset) begin // @[toaxi.scala 77:26]
      raddr <= 32'h0; // @[toaxi.scala 77:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (!(io_dataIO_dc_mode[3])) begin // @[toaxi.scala 101:37]
        if (io_dataIO_dc_mode[2]) begin // @[toaxi.scala 116:43]
          raddr <= io_dataIO_addr; // @[toaxi.scala 129:23]
        end
      end
    end
    if (reset) begin // @[toaxi.scala 78:26]
      rdataEn <= 1'h0; // @[toaxi.scala 78:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_6)) begin // @[Conditional.scala 39:67]
        if (!(_T_8)) begin // @[Conditional.scala 39:67]
          rdataEn <= _GEN_53;
        end
      end
    end
    if (reset) begin // @[toaxi.scala 79:26]
      rdata <= 64'h0; // @[toaxi.scala 79:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_6)) begin // @[Conditional.scala 39:67]
        if (!(_T_8)) begin // @[Conditional.scala 39:67]
          rdata <= _GEN_54;
        end
      end
    end
    if (reset) begin // @[toaxi.scala 81:27]
      pre_addr <= 32'h0; // @[toaxi.scala 81:27]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_dataIO_dc_mode[3]) begin // @[toaxi.scala 101:37]
        pre_addr <= io_dataIO_addr; // @[toaxi.scala 115:26]
      end else if (io_dataIO_dc_mode[2]) begin // @[toaxi.scala 116:43]
        pre_addr <= io_dataIO_addr; // @[toaxi.scala 131:26]
      end
    end
    if (reset) begin // @[toaxi.scala 85:23]
      mode <= 5'h0; // @[toaxi.scala 85:23]
    end else if (_T) begin // @[Conditional.scala 40:58]
      mode <= io_dataIO_dc_mode; // @[toaxi.scala 97:21]
    end
    if (reset) begin // @[toaxi.scala 92:25]
      state <= 3'h0; // @[toaxi.scala 92:25]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_dataIO_dc_mode[3]) begin // @[toaxi.scala 101:37]
        state <= 3'h1; // @[toaxi.scala 102:25]
      end else if (io_dataIO_dc_mode[2]) begin // @[toaxi.scala 116:43]
        state <= 3'h4; // @[toaxi.scala 117:23]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      if (waddrEn & io_outAxi_wa_ready) begin // @[toaxi.scala 136:48]
        state <= 3'h2; // @[toaxi.scala 139:25]
      end
    end else if (_T_8) begin // @[Conditional.scala 39:67]
      state <= _GEN_21;
    end else begin
      state <= _GEN_50;
    end
    if (reset) begin // @[toaxi.scala 208:28]
      out_rdata <= 64'h0; // @[toaxi.scala 208:28]
    end else begin
      out_rdata <= rdata; // @[toaxi.scala 211:15]
    end
    if (reset) begin // @[toaxi.scala 209:28]
      out_valid <= 1'h0; // @[toaxi.scala 209:28]
    end else begin
      out_valid <= state == 3'h6 | state == 3'h3; // @[toaxi.scala 210:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waddrEn = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  waddr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  wsize = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  wdataEn = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  wdata = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  wstrb = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  rsize = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  raddrEn = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  raddr = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  rdataEn = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  rdata = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  pre_addr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  mode = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  state = _RAND_13[2:0];
  _RAND_14 = {2{`RANDOM}};
  out_rdata = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  out_valid = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_CrossBar(
  input         clock,
  input         reset,
  output        io_icAxi_ra_ready,
  input         io_icAxi_ra_valid,
  input  [31:0] io_icAxi_ra_bits_addr,
  output        io_icAxi_rd_valid,
  output [63:0] io_icAxi_rd_bits_data,
  output        io_icAxi_rd_bits_last,
  output        io_flashAxi_wa_ready,
  input         io_flashAxi_wa_valid,
  input  [3:0]  io_flashAxi_wa_bits_id,
  input  [31:0] io_flashAxi_wa_bits_addr,
  input  [7:0]  io_flashAxi_wa_bits_len,
  input  [2:0]  io_flashAxi_wa_bits_size,
  input  [1:0]  io_flashAxi_wa_bits_burst,
  output        io_flashAxi_wd_ready,
  input         io_flashAxi_wd_valid,
  input  [63:0] io_flashAxi_wd_bits_data,
  input  [7:0]  io_flashAxi_wd_bits_strb,
  input         io_flashAxi_wd_bits_last,
  input         io_flashAxi_wr_ready,
  output        io_flashAxi_wr_valid,
  output [3:0]  io_flashAxi_wr_bits_id,
  output [1:0]  io_flashAxi_wr_bits_resp,
  output        io_flashAxi_ra_ready,
  input         io_flashAxi_ra_valid,
  input  [3:0]  io_flashAxi_ra_bits_id,
  input  [31:0] io_flashAxi_ra_bits_addr,
  input  [7:0]  io_flashAxi_ra_bits_len,
  input  [2:0]  io_flashAxi_ra_bits_size,
  input  [1:0]  io_flashAxi_ra_bits_burst,
  input         io_flashAxi_rd_ready,
  output        io_flashAxi_rd_valid,
  output [3:0]  io_flashAxi_rd_bits_id,
  output [63:0] io_flashAxi_rd_bits_data,
  output [1:0]  io_flashAxi_rd_bits_resp,
  output        io_flashAxi_rd_bits_last,
  output        io_memAxi_wa_ready,
  input         io_memAxi_wa_valid,
  input  [31:0] io_memAxi_wa_bits_addr,
  output        io_memAxi_wd_ready,
  input         io_memAxi_wd_valid,
  input  [63:0] io_memAxi_wd_bits_data,
  input         io_memAxi_wd_bits_last,
  output        io_memAxi_ra_ready,
  input         io_memAxi_ra_valid,
  input  [31:0] io_memAxi_ra_bits_addr,
  output        io_memAxi_rd_valid,
  output [63:0] io_memAxi_rd_bits_data,
  output        io_memAxi_rd_bits_last,
  output        io_mmioAxi_wa_ready,
  input         io_mmioAxi_wa_valid,
  input  [3:0]  io_mmioAxi_wa_bits_id,
  input  [31:0] io_mmioAxi_wa_bits_addr,
  input  [7:0]  io_mmioAxi_wa_bits_len,
  input  [2:0]  io_mmioAxi_wa_bits_size,
  input  [1:0]  io_mmioAxi_wa_bits_burst,
  output        io_mmioAxi_wd_ready,
  input         io_mmioAxi_wd_valid,
  input  [63:0] io_mmioAxi_wd_bits_data,
  input  [7:0]  io_mmioAxi_wd_bits_strb,
  input         io_mmioAxi_wd_bits_last,
  input         io_mmioAxi_wr_ready,
  output        io_mmioAxi_wr_valid,
  output [3:0]  io_mmioAxi_wr_bits_id,
  output [1:0]  io_mmioAxi_wr_bits_resp,
  output        io_mmioAxi_ra_ready,
  input         io_mmioAxi_ra_valid,
  input  [3:0]  io_mmioAxi_ra_bits_id,
  input  [31:0] io_mmioAxi_ra_bits_addr,
  input  [7:0]  io_mmioAxi_ra_bits_len,
  input  [2:0]  io_mmioAxi_ra_bits_size,
  input  [1:0]  io_mmioAxi_ra_bits_burst,
  input         io_mmioAxi_rd_ready,
  output        io_mmioAxi_rd_valid,
  output [3:0]  io_mmioAxi_rd_bits_id,
  output [63:0] io_mmioAxi_rd_bits_data,
  output [1:0]  io_mmioAxi_rd_bits_resp,
  output        io_mmioAxi_rd_bits_last,
  input         io_outAxi_wa_ready,
  output        io_outAxi_wa_valid,
  output [3:0]  io_outAxi_wa_bits_id,
  output [31:0] io_outAxi_wa_bits_addr,
  output [7:0]  io_outAxi_wa_bits_len,
  output [2:0]  io_outAxi_wa_bits_size,
  output [1:0]  io_outAxi_wa_bits_burst,
  input         io_outAxi_wd_ready,
  output        io_outAxi_wd_valid,
  output [63:0] io_outAxi_wd_bits_data,
  output [7:0]  io_outAxi_wd_bits_strb,
  output        io_outAxi_wd_bits_last,
  output        io_outAxi_wr_ready,
  input         io_outAxi_wr_valid,
  input  [3:0]  io_outAxi_wr_bits_id,
  input  [1:0]  io_outAxi_wr_bits_resp,
  input         io_outAxi_ra_ready,
  output        io_outAxi_ra_valid,
  output [3:0]  io_outAxi_ra_bits_id,
  output [31:0] io_outAxi_ra_bits_addr,
  output [7:0]  io_outAxi_ra_bits_len,
  output [2:0]  io_outAxi_ra_bits_size,
  output [1:0]  io_outAxi_ra_bits_burst,
  output        io_outAxi_rd_ready,
  input         io_outAxi_rd_valid,
  input  [3:0]  io_outAxi_rd_bits_id,
  input  [63:0] io_outAxi_rd_bits_data,
  input  [1:0]  io_outAxi_rd_bits_resp,
  input         io_outAxi_rd_bits_last,
  input         io_selectMem
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] state; // @[crossbar.scala 20:24]
  reg  selectMem_r; // @[crossbar.scala 22:30]
  wire  memTrans = io_memAxi_ra_valid & io_memAxi_ra_ready | io_memAxi_wa_valid & io_memAxi_wa_ready; // @[crossbar.scala 31:63]
  wire  memDone = io_memAxi_rd_valid & io_memAxi_rd_bits_last | io_memAxi_wd_valid & io_memAxi_wd_ready &
    io_memAxi_wd_bits_last; // @[crossbar.scala 32:88]
  wire  instTrans = io_icAxi_ra_valid & io_icAxi_ra_ready; // @[crossbar.scala 33:40]
  wire  instDone = io_icAxi_rd_valid & io_icAxi_rd_bits_last; // @[crossbar.scala 34:60]
  wire  flashTrans = io_flashAxi_ra_valid & io_flashAxi_ra_ready; // @[crossbar.scala 35:44]
  wire  flashDone = io_flashAxi_rd_valid & io_flashAxi_rd_ready & io_flashAxi_rd_bits_last; // @[crossbar.scala 36:67]
  wire  mmioTrans = io_mmioAxi_ra_valid & io_mmioAxi_ra_ready | io_mmioAxi_wa_valid & io_mmioAxi_wa_ready; // @[crossbar.scala 37:67]
  wire  mmioDone = io_mmioAxi_rd_valid & io_mmioAxi_rd_ready & io_mmioAxi_rd_bits_last | io_mmioAxi_wd_valid &
    io_mmioAxi_wd_ready & io_mmioAxi_wd_bits_last; // @[crossbar.scala 38:93]
  wire  _T = 4'h0 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_0 = io_icAxi_ra_valid ? 4'h2 : state; // @[crossbar.scala 51:42 crossbar.scala 52:23 crossbar.scala 20:24]
  wire [3:0] _GEN_1 = io_flashAxi_ra_valid ? 4'h5 : _GEN_0; // @[crossbar.scala 49:45 crossbar.scala 50:23]
  wire [3:0] _GEN_2 = io_mmioAxi_ra_valid | io_mmioAxi_wa_valid ? 4'h7 : _GEN_1; // @[crossbar.scala 47:67 crossbar.scala 48:23]
  wire  _GEN_5 = io_selectMem | selectMem_r; // @[crossbar.scala 42:31 crossbar.scala 44:29 crossbar.scala 22:30]
  wire  _T_3 = 4'h1 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_6 = memTrans ? 4'h3 : state; // @[crossbar.scala 61:31 crossbar.scala 62:27 crossbar.scala 20:24]
  wire  _GEN_9 = selectMem_r & ~io_selectMem ? 1'h0 : io_outAxi_rd_bits_last; // @[crossbar.scala 56:47 axi.scala 68:23 crossbar.scala 60:27]
  wire [63:0] _GEN_11 = selectMem_r & ~io_selectMem ? 64'h0 : io_outAxi_rd_bits_data; // @[crossbar.scala 56:47 axi.scala 68:23 crossbar.scala 60:27]
  wire  _GEN_13 = selectMem_r & ~io_selectMem ? 1'h0 : io_outAxi_rd_valid; // @[crossbar.scala 56:47 axi.scala 105:18 crossbar.scala 60:27]
  wire  _GEN_14 = selectMem_r & ~io_selectMem ? 1'h0 : 1'h1; // @[crossbar.scala 56:47 axi.scala 87:18 crossbar.scala 60:27]
  wire [1:0] _GEN_15 = selectMem_r & ~io_selectMem ? 2'h0 : 2'h1; // @[crossbar.scala 56:47 axi.scala 41:23 crossbar.scala 60:27]
  wire [2:0] _GEN_16 = selectMem_r & ~io_selectMem ? 3'h0 : 3'h3; // @[crossbar.scala 56:47 axi.scala 41:23 crossbar.scala 60:27]
  wire [7:0] _GEN_17 = selectMem_r & ~io_selectMem ? 8'h0 : 8'h7; // @[crossbar.scala 56:47 axi.scala 41:23 crossbar.scala 60:27]
  wire [31:0] _GEN_18 = selectMem_r & ~io_selectMem ? 32'h0 : io_memAxi_ra_bits_addr; // @[crossbar.scala 56:47 axi.scala 41:23 crossbar.scala 60:27]
  wire  _GEN_20 = selectMem_r & ~io_selectMem ? 1'h0 : io_memAxi_ra_valid; // @[crossbar.scala 56:47 axi.scala 86:18 crossbar.scala 60:27]
  wire  _GEN_21 = selectMem_r & ~io_selectMem ? 1'h0 : io_outAxi_ra_ready; // @[crossbar.scala 56:47 axi.scala 104:18 crossbar.scala 60:27]
  wire  _GEN_26 = selectMem_r & ~io_selectMem ? 1'h0 : io_memAxi_wd_bits_last; // @[crossbar.scala 56:47 axi.scala 50:23 crossbar.scala 60:27]
  wire [7:0] _GEN_27 = selectMem_r & ~io_selectMem ? 8'h0 : 8'hff; // @[crossbar.scala 56:47 axi.scala 50:23 crossbar.scala 60:27]
  wire [63:0] _GEN_28 = selectMem_r & ~io_selectMem ? 64'h0 : io_memAxi_wd_bits_data; // @[crossbar.scala 56:47 axi.scala 50:23 crossbar.scala 60:27]
  wire  _GEN_29 = selectMem_r & ~io_selectMem ? 1'h0 : io_memAxi_wd_valid; // @[crossbar.scala 56:47 axi.scala 84:18 crossbar.scala 60:27]
  wire  _GEN_30 = selectMem_r & ~io_selectMem ? 1'h0 : io_outAxi_wd_ready; // @[crossbar.scala 56:47 axi.scala 102:18 crossbar.scala 60:27]
  wire [31:0] _GEN_34 = selectMem_r & ~io_selectMem ? 32'h0 : io_memAxi_wa_bits_addr; // @[crossbar.scala 56:47 axi.scala 41:23 crossbar.scala 60:27]
  wire  _GEN_36 = selectMem_r & ~io_selectMem ? 1'h0 : io_memAxi_wa_valid; // @[crossbar.scala 56:47 axi.scala 83:18 crossbar.scala 60:27]
  wire  _GEN_37 = selectMem_r & ~io_selectMem ? 1'h0 : io_outAxi_wa_ready; // @[crossbar.scala 56:47 axi.scala 101:18 crossbar.scala 60:27]
  wire  _T_6 = 4'h3 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_38 = memDone ? 4'h0 : state; // @[crossbar.scala 68:26 crossbar.scala 69:23 crossbar.scala 20:24]
  wire  _GEN_39 = memDone ? 1'h0 : selectMem_r; // @[crossbar.scala 68:26 crossbar.scala 70:29 crossbar.scala 22:30]
  wire  _T_7 = 4'h2 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_40 = instTrans ? 4'h4 : state; // @[crossbar.scala 75:28 crossbar.scala 76:23 crossbar.scala 20:24]
  wire  _T_8 = 4'h4 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_41 = instDone ? 4'h0 : state; // @[crossbar.scala 81:27 crossbar.scala 82:23 crossbar.scala 20:24]
  wire  _T_9 = 4'h5 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_42 = flashTrans ? 4'h6 : state; // @[crossbar.scala 87:29 crossbar.scala 88:23 crossbar.scala 20:24]
  wire  _T_10 = 4'h6 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_43 = flashDone ? 4'h0 : state; // @[crossbar.scala 93:28 crossbar.scala 94:23 crossbar.scala 20:24]
  wire  _T_11 = 4'h7 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_44 = mmioTrans ? 4'h8 : state; // @[crossbar.scala 99:28 crossbar.scala 100:23 crossbar.scala 20:24]
  wire  _T_12 = 4'h8 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_45 = mmioDone ? 4'h0 : state; // @[crossbar.scala 105:27 crossbar.scala 106:23 crossbar.scala 20:24]
  wire  _GEN_46 = _T_12 & io_outAxi_rd_bits_last; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 68:23]
  wire [1:0] _GEN_47 = _T_12 ? io_outAxi_rd_bits_resp : 2'h0; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 68:23]
  wire [63:0] _GEN_48 = _T_12 ? io_outAxi_rd_bits_data : 64'h0; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 68:23]
  wire [3:0] _GEN_49 = _T_12 ? io_outAxi_rd_bits_id : 4'h0; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 68:23]
  wire  _GEN_50 = _T_12 & io_outAxi_rd_valid; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 105:18]
  wire  _GEN_51 = _T_12 & io_mmioAxi_rd_ready; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 87:18]
  wire [1:0] _GEN_52 = _T_12 ? io_mmioAxi_ra_bits_burst : 2'h0; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 41:23]
  wire [2:0] _GEN_53 = _T_12 ? io_mmioAxi_ra_bits_size : 3'h0; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 41:23]
  wire [7:0] _GEN_54 = _T_12 ? io_mmioAxi_ra_bits_len : 8'h0; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 41:23]
  wire [31:0] _GEN_55 = _T_12 ? io_mmioAxi_ra_bits_addr : 32'h0; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 41:23]
  wire [3:0] _GEN_56 = _T_12 ? io_mmioAxi_ra_bits_id : 4'h0; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 41:23]
  wire  _GEN_57 = _T_12 & io_mmioAxi_ra_valid; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 86:18]
  wire  _GEN_58 = _T_12 & io_outAxi_ra_ready; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 104:18]
  wire [1:0] _GEN_59 = _T_12 ? io_outAxi_wr_bits_resp : 2'h0; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 58:23]
  wire [3:0] _GEN_60 = _T_12 ? io_outAxi_wr_bits_id : 4'h0; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 58:23]
  wire  _GEN_61 = _T_12 & io_outAxi_wr_valid; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 103:18]
  wire  _GEN_62 = _T_12 ? io_mmioAxi_wr_ready : 1'h1; // @[Conditional.scala 39:67 crossbar.scala 104:23 crossbar.scala 29:24]
  wire  _GEN_63 = _T_12 & io_mmioAxi_wd_bits_last; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 50:23]
  wire [7:0] _GEN_64 = _T_12 ? io_mmioAxi_wd_bits_strb : 8'h0; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 50:23]
  wire [63:0] _GEN_65 = _T_12 ? io_mmioAxi_wd_bits_data : 64'h0; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 50:23]
  wire  _GEN_66 = _T_12 & io_mmioAxi_wd_valid; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 84:18]
  wire  _GEN_67 = _T_12 & io_outAxi_wd_ready; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 102:18]
  wire [1:0] _GEN_68 = _T_12 ? io_mmioAxi_wa_bits_burst : 2'h0; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 41:23]
  wire [2:0] _GEN_69 = _T_12 ? io_mmioAxi_wa_bits_size : 3'h0; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 41:23]
  wire [7:0] _GEN_70 = _T_12 ? io_mmioAxi_wa_bits_len : 8'h0; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 41:23]
  wire [31:0] _GEN_71 = _T_12 ? io_mmioAxi_wa_bits_addr : 32'h0; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 41:23]
  wire [3:0] _GEN_72 = _T_12 ? io_mmioAxi_wa_bits_id : 4'h0; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 41:23]
  wire  _GEN_73 = _T_12 & io_mmioAxi_wa_valid; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 83:18]
  wire  _GEN_74 = _T_12 & io_outAxi_wa_ready; // @[Conditional.scala 39:67 crossbar.scala 104:23 axi.scala 101:18]
  wire [3:0] _GEN_75 = _T_12 ? _GEN_45 : state; // @[Conditional.scala 39:67 crossbar.scala 20:24]
  wire  _GEN_76 = _T_11 ? io_outAxi_rd_bits_last : _GEN_46; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [1:0] _GEN_77 = _T_11 ? io_outAxi_rd_bits_resp : _GEN_47; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [63:0] _GEN_78 = _T_11 ? io_outAxi_rd_bits_data : _GEN_48; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [3:0] _GEN_79 = _T_11 ? io_outAxi_rd_bits_id : _GEN_49; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire  _GEN_80 = _T_11 ? io_outAxi_rd_valid : _GEN_50; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire  _GEN_81 = _T_11 ? io_mmioAxi_rd_ready : _GEN_51; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [1:0] _GEN_82 = _T_11 ? io_mmioAxi_ra_bits_burst : _GEN_52; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [2:0] _GEN_83 = _T_11 ? io_mmioAxi_ra_bits_size : _GEN_53; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [7:0] _GEN_84 = _T_11 ? io_mmioAxi_ra_bits_len : _GEN_54; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [31:0] _GEN_85 = _T_11 ? io_mmioAxi_ra_bits_addr : _GEN_55; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [3:0] _GEN_86 = _T_11 ? io_mmioAxi_ra_bits_id : _GEN_56; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire  _GEN_87 = _T_11 ? io_mmioAxi_ra_valid : _GEN_57; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire  _GEN_88 = _T_11 ? io_outAxi_ra_ready : _GEN_58; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [1:0] _GEN_89 = _T_11 ? io_outAxi_wr_bits_resp : _GEN_59; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [3:0] _GEN_90 = _T_11 ? io_outAxi_wr_bits_id : _GEN_60; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire  _GEN_91 = _T_11 ? io_outAxi_wr_valid : _GEN_61; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire  _GEN_92 = _T_11 ? io_mmioAxi_wr_ready : _GEN_62; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire  _GEN_93 = _T_11 ? io_mmioAxi_wd_bits_last : _GEN_63; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [7:0] _GEN_94 = _T_11 ? io_mmioAxi_wd_bits_strb : _GEN_64; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [63:0] _GEN_95 = _T_11 ? io_mmioAxi_wd_bits_data : _GEN_65; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire  _GEN_96 = _T_11 ? io_mmioAxi_wd_valid : _GEN_66; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire  _GEN_97 = _T_11 ? io_outAxi_wd_ready : _GEN_67; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [1:0] _GEN_98 = _T_11 ? io_mmioAxi_wa_bits_burst : _GEN_68; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [2:0] _GEN_99 = _T_11 ? io_mmioAxi_wa_bits_size : _GEN_69; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [7:0] _GEN_100 = _T_11 ? io_mmioAxi_wa_bits_len : _GEN_70; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [31:0] _GEN_101 = _T_11 ? io_mmioAxi_wa_bits_addr : _GEN_71; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [3:0] _GEN_102 = _T_11 ? io_mmioAxi_wa_bits_id : _GEN_72; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire  _GEN_103 = _T_11 ? io_mmioAxi_wa_valid : _GEN_73; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire  _GEN_104 = _T_11 ? io_outAxi_wa_ready : _GEN_74; // @[Conditional.scala 39:67 crossbar.scala 98:23]
  wire [3:0] _GEN_105 = _T_11 ? _GEN_44 : _GEN_75; // @[Conditional.scala 39:67]
  wire  _GEN_106 = _T_10 & io_outAxi_rd_bits_last; // @[Conditional.scala 39:67 crossbar.scala 92:23 axi.scala 68:23]
  wire [1:0] _GEN_107 = _T_10 ? io_outAxi_rd_bits_resp : 2'h0; // @[Conditional.scala 39:67 crossbar.scala 92:23 axi.scala 68:23]
  wire [63:0] _GEN_108 = _T_10 ? io_outAxi_rd_bits_data : 64'h0; // @[Conditional.scala 39:67 crossbar.scala 92:23 axi.scala 68:23]
  wire [3:0] _GEN_109 = _T_10 ? io_outAxi_rd_bits_id : 4'h0; // @[Conditional.scala 39:67 crossbar.scala 92:23 axi.scala 68:23]
  wire  _GEN_110 = _T_10 & io_outAxi_rd_valid; // @[Conditional.scala 39:67 crossbar.scala 92:23 axi.scala 105:18]
  wire  _GEN_111 = _T_10 ? io_flashAxi_rd_ready : _GEN_81; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire [1:0] _GEN_112 = _T_10 ? io_flashAxi_ra_bits_burst : _GEN_82; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire [2:0] _GEN_113 = _T_10 ? io_flashAxi_ra_bits_size : _GEN_83; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire [7:0] _GEN_114 = _T_10 ? io_flashAxi_ra_bits_len : _GEN_84; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire [31:0] _GEN_115 = _T_10 ? io_flashAxi_ra_bits_addr : _GEN_85; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire [3:0] _GEN_116 = _T_10 ? io_flashAxi_ra_bits_id : _GEN_86; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire  _GEN_117 = _T_10 ? io_flashAxi_ra_valid : _GEN_87; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire  _GEN_118 = _T_10 & io_outAxi_ra_ready; // @[Conditional.scala 39:67 crossbar.scala 92:23 axi.scala 104:18]
  wire [1:0] _GEN_119 = _T_10 ? io_outAxi_wr_bits_resp : 2'h0; // @[Conditional.scala 39:67 crossbar.scala 92:23 axi.scala 58:23]
  wire [3:0] _GEN_120 = _T_10 ? io_outAxi_wr_bits_id : 4'h0; // @[Conditional.scala 39:67 crossbar.scala 92:23 axi.scala 58:23]
  wire  _GEN_121 = _T_10 & io_outAxi_wr_valid; // @[Conditional.scala 39:67 crossbar.scala 92:23 axi.scala 103:18]
  wire  _GEN_122 = _T_10 ? io_flashAxi_wr_ready : _GEN_92; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire  _GEN_123 = _T_10 ? io_flashAxi_wd_bits_last : _GEN_93; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire [7:0] _GEN_124 = _T_10 ? io_flashAxi_wd_bits_strb : _GEN_94; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire [63:0] _GEN_125 = _T_10 ? io_flashAxi_wd_bits_data : _GEN_95; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire  _GEN_126 = _T_10 ? io_flashAxi_wd_valid : _GEN_96; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire  _GEN_127 = _T_10 & io_outAxi_wd_ready; // @[Conditional.scala 39:67 crossbar.scala 92:23 axi.scala 102:18]
  wire [1:0] _GEN_128 = _T_10 ? io_flashAxi_wa_bits_burst : _GEN_98; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire [2:0] _GEN_129 = _T_10 ? io_flashAxi_wa_bits_size : _GEN_99; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire [7:0] _GEN_130 = _T_10 ? io_flashAxi_wa_bits_len : _GEN_100; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire [31:0] _GEN_131 = _T_10 ? io_flashAxi_wa_bits_addr : _GEN_101; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire [3:0] _GEN_132 = _T_10 ? io_flashAxi_wa_bits_id : _GEN_102; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire  _GEN_133 = _T_10 ? io_flashAxi_wa_valid : _GEN_103; // @[Conditional.scala 39:67 crossbar.scala 92:23]
  wire  _GEN_134 = _T_10 & io_outAxi_wa_ready; // @[Conditional.scala 39:67 crossbar.scala 92:23 axi.scala 101:18]
  wire [3:0] _GEN_135 = _T_10 ? _GEN_43 : _GEN_105; // @[Conditional.scala 39:67]
  wire  _GEN_136 = _T_10 ? 1'h0 : _GEN_76; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [1:0] _GEN_137 = _T_10 ? 2'h0 : _GEN_77; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [63:0] _GEN_138 = _T_10 ? 64'h0 : _GEN_78; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [3:0] _GEN_139 = _T_10 ? 4'h0 : _GEN_79; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire  _GEN_140 = _T_10 ? 1'h0 : _GEN_80; // @[Conditional.scala 39:67 axi.scala 105:18]
  wire  _GEN_141 = _T_10 ? 1'h0 : _GEN_88; // @[Conditional.scala 39:67 axi.scala 104:18]
  wire [1:0] _GEN_142 = _T_10 ? 2'h0 : _GEN_89; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire [3:0] _GEN_143 = _T_10 ? 4'h0 : _GEN_90; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire  _GEN_144 = _T_10 ? 1'h0 : _GEN_91; // @[Conditional.scala 39:67 axi.scala 103:18]
  wire  _GEN_145 = _T_10 ? 1'h0 : _GEN_97; // @[Conditional.scala 39:67 axi.scala 102:18]
  wire  _GEN_146 = _T_10 ? 1'h0 : _GEN_104; // @[Conditional.scala 39:67 axi.scala 101:18]
  wire  _GEN_147 = _T_9 ? io_outAxi_rd_bits_last : _GEN_106; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [1:0] _GEN_148 = _T_9 ? io_outAxi_rd_bits_resp : _GEN_107; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [63:0] _GEN_149 = _T_9 ? io_outAxi_rd_bits_data : _GEN_108; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [3:0] _GEN_150 = _T_9 ? io_outAxi_rd_bits_id : _GEN_109; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire  _GEN_151 = _T_9 ? io_outAxi_rd_valid : _GEN_110; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire  _GEN_152 = _T_9 ? io_flashAxi_rd_ready : _GEN_111; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [1:0] _GEN_153 = _T_9 ? io_flashAxi_ra_bits_burst : _GEN_112; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [2:0] _GEN_154 = _T_9 ? io_flashAxi_ra_bits_size : _GEN_113; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [7:0] _GEN_155 = _T_9 ? io_flashAxi_ra_bits_len : _GEN_114; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [31:0] _GEN_156 = _T_9 ? io_flashAxi_ra_bits_addr : _GEN_115; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [3:0] _GEN_157 = _T_9 ? io_flashAxi_ra_bits_id : _GEN_116; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire  _GEN_158 = _T_9 ? io_flashAxi_ra_valid : _GEN_117; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire  _GEN_159 = _T_9 ? io_outAxi_ra_ready : _GEN_118; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [1:0] _GEN_160 = _T_9 ? io_outAxi_wr_bits_resp : _GEN_119; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [3:0] _GEN_161 = _T_9 ? io_outAxi_wr_bits_id : _GEN_120; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire  _GEN_162 = _T_9 ? io_outAxi_wr_valid : _GEN_121; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire  _GEN_163 = _T_9 ? io_flashAxi_wr_ready : _GEN_122; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire  _GEN_164 = _T_9 ? io_flashAxi_wd_bits_last : _GEN_123; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [7:0] _GEN_165 = _T_9 ? io_flashAxi_wd_bits_strb : _GEN_124; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [63:0] _GEN_166 = _T_9 ? io_flashAxi_wd_bits_data : _GEN_125; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire  _GEN_167 = _T_9 ? io_flashAxi_wd_valid : _GEN_126; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire  _GEN_168 = _T_9 ? io_outAxi_wd_ready : _GEN_127; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [1:0] _GEN_169 = _T_9 ? io_flashAxi_wa_bits_burst : _GEN_128; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [2:0] _GEN_170 = _T_9 ? io_flashAxi_wa_bits_size : _GEN_129; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [7:0] _GEN_171 = _T_9 ? io_flashAxi_wa_bits_len : _GEN_130; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [31:0] _GEN_172 = _T_9 ? io_flashAxi_wa_bits_addr : _GEN_131; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [3:0] _GEN_173 = _T_9 ? io_flashAxi_wa_bits_id : _GEN_132; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire  _GEN_174 = _T_9 ? io_flashAxi_wa_valid : _GEN_133; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire  _GEN_175 = _T_9 ? io_outAxi_wa_ready : _GEN_134; // @[Conditional.scala 39:67 crossbar.scala 86:23]
  wire [3:0] _GEN_176 = _T_9 ? _GEN_42 : _GEN_135; // @[Conditional.scala 39:67]
  wire  _GEN_177 = _T_9 ? 1'h0 : _GEN_136; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [1:0] _GEN_178 = _T_9 ? 2'h0 : _GEN_137; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [63:0] _GEN_179 = _T_9 ? 64'h0 : _GEN_138; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [3:0] _GEN_180 = _T_9 ? 4'h0 : _GEN_139; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire  _GEN_181 = _T_9 ? 1'h0 : _GEN_140; // @[Conditional.scala 39:67 axi.scala 105:18]
  wire  _GEN_182 = _T_9 ? 1'h0 : _GEN_141; // @[Conditional.scala 39:67 axi.scala 104:18]
  wire [1:0] _GEN_183 = _T_9 ? 2'h0 : _GEN_142; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire [3:0] _GEN_184 = _T_9 ? 4'h0 : _GEN_143; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire  _GEN_185 = _T_9 ? 1'h0 : _GEN_144; // @[Conditional.scala 39:67 axi.scala 103:18]
  wire  _GEN_186 = _T_9 ? 1'h0 : _GEN_145; // @[Conditional.scala 39:67 axi.scala 102:18]
  wire  _GEN_187 = _T_9 ? 1'h0 : _GEN_146; // @[Conditional.scala 39:67 axi.scala 101:18]
  wire  _GEN_188 = _T_8 & io_outAxi_rd_bits_last; // @[Conditional.scala 39:67 crossbar.scala 80:23 axi.scala 68:23]
  wire [63:0] _GEN_190 = _T_8 ? io_outAxi_rd_bits_data : 64'h0; // @[Conditional.scala 39:67 crossbar.scala 80:23 axi.scala 68:23]
  wire  _GEN_192 = _T_8 & io_outAxi_rd_valid; // @[Conditional.scala 39:67 crossbar.scala 80:23 axi.scala 105:18]
  wire  _GEN_193 = _T_8 | _GEN_152; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire [1:0] _GEN_194 = _T_8 ? 2'h1 : _GEN_153; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire [2:0] _GEN_195 = _T_8 ? 3'h3 : _GEN_154; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire [7:0] _GEN_196 = _T_8 ? 8'h7 : _GEN_155; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire [31:0] _GEN_197 = _T_8 ? io_icAxi_ra_bits_addr : _GEN_156; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire [3:0] _GEN_198 = _T_8 ? 4'h0 : _GEN_157; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire  _GEN_199 = _T_8 ? io_icAxi_ra_valid : _GEN_158; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire  _GEN_200 = _T_8 & io_outAxi_ra_ready; // @[Conditional.scala 39:67 crossbar.scala 80:23 axi.scala 104:18]
  wire  _GEN_204 = _T_8 | _GEN_163; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire  _GEN_205 = _T_8 ? 1'h0 : _GEN_164; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire [7:0] _GEN_206 = _T_8 ? 8'h0 : _GEN_165; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire [63:0] _GEN_207 = _T_8 ? 64'h0 : _GEN_166; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire  _GEN_208 = _T_8 ? 1'h0 : _GEN_167; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire [1:0] _GEN_210 = _T_8 ? 2'h0 : _GEN_169; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire [2:0] _GEN_211 = _T_8 ? 3'h0 : _GEN_170; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire [7:0] _GEN_212 = _T_8 ? 8'h0 : _GEN_171; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire [31:0] _GEN_213 = _T_8 ? 32'h0 : _GEN_172; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire [3:0] _GEN_214 = _T_8 ? 4'h0 : _GEN_173; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire  _GEN_215 = _T_8 ? 1'h0 : _GEN_174; // @[Conditional.scala 39:67 crossbar.scala 80:23]
  wire [3:0] _GEN_217 = _T_8 ? _GEN_41 : _GEN_176; // @[Conditional.scala 39:67]
  wire  _GEN_218 = _T_8 ? 1'h0 : _GEN_147; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [1:0] _GEN_219 = _T_8 ? 2'h0 : _GEN_148; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [63:0] _GEN_220 = _T_8 ? 64'h0 : _GEN_149; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [3:0] _GEN_221 = _T_8 ? 4'h0 : _GEN_150; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire  _GEN_222 = _T_8 ? 1'h0 : _GEN_151; // @[Conditional.scala 39:67 axi.scala 105:18]
  wire  _GEN_223 = _T_8 ? 1'h0 : _GEN_159; // @[Conditional.scala 39:67 axi.scala 104:18]
  wire [1:0] _GEN_224 = _T_8 ? 2'h0 : _GEN_160; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire [3:0] _GEN_225 = _T_8 ? 4'h0 : _GEN_161; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire  _GEN_226 = _T_8 ? 1'h0 : _GEN_162; // @[Conditional.scala 39:67 axi.scala 103:18]
  wire  _GEN_227 = _T_8 ? 1'h0 : _GEN_168; // @[Conditional.scala 39:67 axi.scala 102:18]
  wire  _GEN_228 = _T_8 ? 1'h0 : _GEN_175; // @[Conditional.scala 39:67 axi.scala 101:18]
  wire  _GEN_229 = _T_8 ? 1'h0 : _GEN_177; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [1:0] _GEN_230 = _T_8 ? 2'h0 : _GEN_178; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [63:0] _GEN_231 = _T_8 ? 64'h0 : _GEN_179; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [3:0] _GEN_232 = _T_8 ? 4'h0 : _GEN_180; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire  _GEN_233 = _T_8 ? 1'h0 : _GEN_181; // @[Conditional.scala 39:67 axi.scala 105:18]
  wire  _GEN_234 = _T_8 ? 1'h0 : _GEN_182; // @[Conditional.scala 39:67 axi.scala 104:18]
  wire [1:0] _GEN_235 = _T_8 ? 2'h0 : _GEN_183; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire [3:0] _GEN_236 = _T_8 ? 4'h0 : _GEN_184; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire  _GEN_237 = _T_8 ? 1'h0 : _GEN_185; // @[Conditional.scala 39:67 axi.scala 103:18]
  wire  _GEN_238 = _T_8 ? 1'h0 : _GEN_186; // @[Conditional.scala 39:67 axi.scala 102:18]
  wire  _GEN_239 = _T_8 ? 1'h0 : _GEN_187; // @[Conditional.scala 39:67 axi.scala 101:18]
  wire  _GEN_240 = _T_7 ? io_outAxi_rd_bits_last : _GEN_188; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire [63:0] _GEN_242 = _T_7 ? io_outAxi_rd_bits_data : _GEN_190; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire  _GEN_244 = _T_7 ? io_outAxi_rd_valid : _GEN_192; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire  _GEN_245 = _T_7 | _GEN_193; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire [1:0] _GEN_246 = _T_7 ? 2'h1 : _GEN_194; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire [2:0] _GEN_247 = _T_7 ? 3'h3 : _GEN_195; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire [7:0] _GEN_248 = _T_7 ? 8'h7 : _GEN_196; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire [31:0] _GEN_249 = _T_7 ? io_icAxi_ra_bits_addr : _GEN_197; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire [3:0] _GEN_250 = _T_7 ? 4'h0 : _GEN_198; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire  _GEN_251 = _T_7 ? io_icAxi_ra_valid : _GEN_199; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire  _GEN_252 = _T_7 ? io_outAxi_ra_ready : _GEN_200; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire  _GEN_256 = _T_7 | _GEN_204; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire  _GEN_257 = _T_7 ? 1'h0 : _GEN_205; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire [7:0] _GEN_258 = _T_7 ? 8'h0 : _GEN_206; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire [63:0] _GEN_259 = _T_7 ? 64'h0 : _GEN_207; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire  _GEN_260 = _T_7 ? 1'h0 : _GEN_208; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire [1:0] _GEN_262 = _T_7 ? 2'h0 : _GEN_210; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire [2:0] _GEN_263 = _T_7 ? 3'h0 : _GEN_211; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire [7:0] _GEN_264 = _T_7 ? 8'h0 : _GEN_212; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire [31:0] _GEN_265 = _T_7 ? 32'h0 : _GEN_213; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire [3:0] _GEN_266 = _T_7 ? 4'h0 : _GEN_214; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire  _GEN_267 = _T_7 ? 1'h0 : _GEN_215; // @[Conditional.scala 39:67 crossbar.scala 74:23]
  wire [3:0] _GEN_269 = _T_7 ? _GEN_40 : _GEN_217; // @[Conditional.scala 39:67]
  wire  _GEN_270 = _T_7 ? 1'h0 : _GEN_218; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [1:0] _GEN_271 = _T_7 ? 2'h0 : _GEN_219; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [63:0] _GEN_272 = _T_7 ? 64'h0 : _GEN_220; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [3:0] _GEN_273 = _T_7 ? 4'h0 : _GEN_221; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire  _GEN_274 = _T_7 ? 1'h0 : _GEN_222; // @[Conditional.scala 39:67 axi.scala 105:18]
  wire  _GEN_275 = _T_7 ? 1'h0 : _GEN_223; // @[Conditional.scala 39:67 axi.scala 104:18]
  wire [1:0] _GEN_276 = _T_7 ? 2'h0 : _GEN_224; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire [3:0] _GEN_277 = _T_7 ? 4'h0 : _GEN_225; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire  _GEN_278 = _T_7 ? 1'h0 : _GEN_226; // @[Conditional.scala 39:67 axi.scala 103:18]
  wire  _GEN_279 = _T_7 ? 1'h0 : _GEN_227; // @[Conditional.scala 39:67 axi.scala 102:18]
  wire  _GEN_280 = _T_7 ? 1'h0 : _GEN_228; // @[Conditional.scala 39:67 axi.scala 101:18]
  wire  _GEN_281 = _T_7 ? 1'h0 : _GEN_229; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [1:0] _GEN_282 = _T_7 ? 2'h0 : _GEN_230; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [63:0] _GEN_283 = _T_7 ? 64'h0 : _GEN_231; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [3:0] _GEN_284 = _T_7 ? 4'h0 : _GEN_232; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire  _GEN_285 = _T_7 ? 1'h0 : _GEN_233; // @[Conditional.scala 39:67 axi.scala 105:18]
  wire  _GEN_286 = _T_7 ? 1'h0 : _GEN_234; // @[Conditional.scala 39:67 axi.scala 104:18]
  wire [1:0] _GEN_287 = _T_7 ? 2'h0 : _GEN_235; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire [3:0] _GEN_288 = _T_7 ? 4'h0 : _GEN_236; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire  _GEN_289 = _T_7 ? 1'h0 : _GEN_237; // @[Conditional.scala 39:67 axi.scala 103:18]
  wire  _GEN_290 = _T_7 ? 1'h0 : _GEN_238; // @[Conditional.scala 39:67 axi.scala 102:18]
  wire  _GEN_291 = _T_7 ? 1'h0 : _GEN_239; // @[Conditional.scala 39:67 axi.scala 101:18]
  wire  _GEN_292 = _T_6 & io_outAxi_rd_bits_last; // @[Conditional.scala 39:67 crossbar.scala 67:23 axi.scala 68:23]
  wire [63:0] _GEN_294 = _T_6 ? io_outAxi_rd_bits_data : 64'h0; // @[Conditional.scala 39:67 crossbar.scala 67:23 axi.scala 68:23]
  wire  _GEN_296 = _T_6 & io_outAxi_rd_valid; // @[Conditional.scala 39:67 crossbar.scala 67:23 axi.scala 105:18]
  wire  _GEN_297 = _T_6 | _GEN_245; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire [1:0] _GEN_298 = _T_6 ? 2'h1 : _GEN_246; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire [2:0] _GEN_299 = _T_6 ? 3'h3 : _GEN_247; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire [7:0] _GEN_300 = _T_6 ? 8'h7 : _GEN_248; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire [31:0] _GEN_301 = _T_6 ? io_memAxi_ra_bits_addr : _GEN_249; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire [3:0] _GEN_302 = _T_6 ? 4'h0 : _GEN_250; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire  _GEN_303 = _T_6 ? io_memAxi_ra_valid : _GEN_251; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire  _GEN_304 = _T_6 & io_outAxi_ra_ready; // @[Conditional.scala 39:67 crossbar.scala 67:23 axi.scala 104:18]
  wire  _GEN_308 = _T_6 | _GEN_256; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire  _GEN_309 = _T_6 ? io_memAxi_wd_bits_last : _GEN_257; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire [7:0] _GEN_310 = _T_6 ? 8'hff : _GEN_258; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire [63:0] _GEN_311 = _T_6 ? io_memAxi_wd_bits_data : _GEN_259; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire  _GEN_312 = _T_6 ? io_memAxi_wd_valid : _GEN_260; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire  _GEN_313 = _T_6 & io_outAxi_wd_ready; // @[Conditional.scala 39:67 crossbar.scala 67:23 axi.scala 102:18]
  wire [1:0] _GEN_314 = _T_6 ? 2'h1 : _GEN_262; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire [2:0] _GEN_315 = _T_6 ? 3'h3 : _GEN_263; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire [7:0] _GEN_316 = _T_6 ? 8'h7 : _GEN_264; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire [31:0] _GEN_317 = _T_6 ? io_memAxi_wa_bits_addr : _GEN_265; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire [3:0] _GEN_318 = _T_6 ? 4'h0 : _GEN_266; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire  _GEN_319 = _T_6 ? io_memAxi_wa_valid : _GEN_267; // @[Conditional.scala 39:67 crossbar.scala 67:23]
  wire  _GEN_320 = _T_6 & io_outAxi_wa_ready; // @[Conditional.scala 39:67 crossbar.scala 67:23 axi.scala 101:18]
  wire  _GEN_323 = _T_6 ? 1'h0 : _GEN_240; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [63:0] _GEN_325 = _T_6 ? 64'h0 : _GEN_242; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire  _GEN_327 = _T_6 ? 1'h0 : _GEN_244; // @[Conditional.scala 39:67 axi.scala 105:18]
  wire  _GEN_328 = _T_6 ? 1'h0 : _GEN_252; // @[Conditional.scala 39:67 axi.scala 104:18]
  wire  _GEN_334 = _T_6 ? 1'h0 : _GEN_270; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [1:0] _GEN_335 = _T_6 ? 2'h0 : _GEN_271; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [63:0] _GEN_336 = _T_6 ? 64'h0 : _GEN_272; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [3:0] _GEN_337 = _T_6 ? 4'h0 : _GEN_273; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire  _GEN_338 = _T_6 ? 1'h0 : _GEN_274; // @[Conditional.scala 39:67 axi.scala 105:18]
  wire  _GEN_339 = _T_6 ? 1'h0 : _GEN_275; // @[Conditional.scala 39:67 axi.scala 104:18]
  wire [1:0] _GEN_340 = _T_6 ? 2'h0 : _GEN_276; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire [3:0] _GEN_341 = _T_6 ? 4'h0 : _GEN_277; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire  _GEN_342 = _T_6 ? 1'h0 : _GEN_278; // @[Conditional.scala 39:67 axi.scala 103:18]
  wire  _GEN_343 = _T_6 ? 1'h0 : _GEN_279; // @[Conditional.scala 39:67 axi.scala 102:18]
  wire  _GEN_344 = _T_6 ? 1'h0 : _GEN_280; // @[Conditional.scala 39:67 axi.scala 101:18]
  wire  _GEN_345 = _T_6 ? 1'h0 : _GEN_281; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [1:0] _GEN_346 = _T_6 ? 2'h0 : _GEN_282; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [63:0] _GEN_347 = _T_6 ? 64'h0 : _GEN_283; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [3:0] _GEN_348 = _T_6 ? 4'h0 : _GEN_284; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire  _GEN_349 = _T_6 ? 1'h0 : _GEN_285; // @[Conditional.scala 39:67 axi.scala 105:18]
  wire  _GEN_350 = _T_6 ? 1'h0 : _GEN_286; // @[Conditional.scala 39:67 axi.scala 104:18]
  wire [1:0] _GEN_351 = _T_6 ? 2'h0 : _GEN_287; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire [3:0] _GEN_352 = _T_6 ? 4'h0 : _GEN_288; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire  _GEN_353 = _T_6 ? 1'h0 : _GEN_289; // @[Conditional.scala 39:67 axi.scala 103:18]
  wire  _GEN_354 = _T_6 ? 1'h0 : _GEN_290; // @[Conditional.scala 39:67 axi.scala 102:18]
  wire  _GEN_355 = _T_6 ? 1'h0 : _GEN_291; // @[Conditional.scala 39:67 axi.scala 101:18]
  wire  _GEN_358 = _T_3 ? _GEN_9 : _GEN_292; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_360 = _T_3 ? _GEN_11 : _GEN_294; // @[Conditional.scala 39:67]
  wire  _GEN_362 = _T_3 ? _GEN_13 : _GEN_296; // @[Conditional.scala 39:67]
  wire  _GEN_363 = _T_3 ? _GEN_14 : _GEN_297; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_364 = _T_3 ? _GEN_15 : _GEN_298; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_365 = _T_3 ? _GEN_16 : _GEN_299; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_366 = _T_3 ? _GEN_17 : _GEN_300; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_367 = _T_3 ? _GEN_18 : _GEN_301; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_368 = _T_3 ? 4'h0 : _GEN_302; // @[Conditional.scala 39:67]
  wire  _GEN_369 = _T_3 ? _GEN_20 : _GEN_303; // @[Conditional.scala 39:67]
  wire  _GEN_370 = _T_3 ? _GEN_21 : _GEN_304; // @[Conditional.scala 39:67]
  wire  _GEN_374 = _T_3 | _GEN_308; // @[Conditional.scala 39:67]
  wire  _GEN_375 = _T_3 ? _GEN_26 : _GEN_309; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_376 = _T_3 ? _GEN_27 : _GEN_310; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_377 = _T_3 ? _GEN_28 : _GEN_311; // @[Conditional.scala 39:67]
  wire  _GEN_378 = _T_3 ? _GEN_29 : _GEN_312; // @[Conditional.scala 39:67]
  wire  _GEN_379 = _T_3 ? _GEN_30 : _GEN_313; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_380 = _T_3 ? _GEN_15 : _GEN_314; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_381 = _T_3 ? _GEN_16 : _GEN_315; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_382 = _T_3 ? _GEN_17 : _GEN_316; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_383 = _T_3 ? _GEN_34 : _GEN_317; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_384 = _T_3 ? 4'h0 : _GEN_318; // @[Conditional.scala 39:67]
  wire  _GEN_385 = _T_3 ? _GEN_36 : _GEN_319; // @[Conditional.scala 39:67]
  wire  _GEN_386 = _T_3 ? _GEN_37 : _GEN_320; // @[Conditional.scala 39:67]
  wire  _GEN_387 = _T_3 ? 1'h0 : _GEN_323; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [63:0] _GEN_389 = _T_3 ? 64'h0 : _GEN_325; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire  _GEN_391 = _T_3 ? 1'h0 : _GEN_327; // @[Conditional.scala 39:67 axi.scala 105:18]
  wire  _GEN_392 = _T_3 ? 1'h0 : _GEN_328; // @[Conditional.scala 39:67 axi.scala 104:18]
  wire  _GEN_398 = _T_3 ? 1'h0 : _GEN_334; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [1:0] _GEN_399 = _T_3 ? 2'h0 : _GEN_335; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [63:0] _GEN_400 = _T_3 ? 64'h0 : _GEN_336; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [3:0] _GEN_401 = _T_3 ? 4'h0 : _GEN_337; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire  _GEN_402 = _T_3 ? 1'h0 : _GEN_338; // @[Conditional.scala 39:67 axi.scala 105:18]
  wire  _GEN_403 = _T_3 ? 1'h0 : _GEN_339; // @[Conditional.scala 39:67 axi.scala 104:18]
  wire [1:0] _GEN_404 = _T_3 ? 2'h0 : _GEN_340; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire [3:0] _GEN_405 = _T_3 ? 4'h0 : _GEN_341; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire  _GEN_406 = _T_3 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 axi.scala 103:18]
  wire  _GEN_407 = _T_3 ? 1'h0 : _GEN_343; // @[Conditional.scala 39:67 axi.scala 102:18]
  wire  _GEN_408 = _T_3 ? 1'h0 : _GEN_344; // @[Conditional.scala 39:67 axi.scala 101:18]
  wire  _GEN_409 = _T_3 ? 1'h0 : _GEN_345; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [1:0] _GEN_410 = _T_3 ? 2'h0 : _GEN_346; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [63:0] _GEN_411 = _T_3 ? 64'h0 : _GEN_347; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire [3:0] _GEN_412 = _T_3 ? 4'h0 : _GEN_348; // @[Conditional.scala 39:67 axi.scala 68:23]
  wire  _GEN_413 = _T_3 ? 1'h0 : _GEN_349; // @[Conditional.scala 39:67 axi.scala 105:18]
  wire  _GEN_414 = _T_3 ? 1'h0 : _GEN_350; // @[Conditional.scala 39:67 axi.scala 104:18]
  wire [1:0] _GEN_415 = _T_3 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire [3:0] _GEN_416 = _T_3 ? 4'h0 : _GEN_352; // @[Conditional.scala 39:67 axi.scala 58:23]
  wire  _GEN_417 = _T_3 ? 1'h0 : _GEN_353; // @[Conditional.scala 39:67 axi.scala 103:18]
  wire  _GEN_418 = _T_3 ? 1'h0 : _GEN_354; // @[Conditional.scala 39:67 axi.scala 102:18]
  wire  _GEN_419 = _T_3 ? 1'h0 : _GEN_355; // @[Conditional.scala 39:67 axi.scala 101:18]
  assign io_icAxi_ra_ready = _T ? 1'h0 : _GEN_392; // @[Conditional.scala 40:58 axi.scala 104:18]
  assign io_icAxi_rd_valid = _T ? 1'h0 : _GEN_391; // @[Conditional.scala 40:58 axi.scala 105:18]
  assign io_icAxi_rd_bits_data = _T ? 64'h0 : _GEN_389; // @[Conditional.scala 40:58 axi.scala 68:23]
  assign io_icAxi_rd_bits_last = _T ? 1'h0 : _GEN_387; // @[Conditional.scala 40:58 axi.scala 68:23]
  assign io_flashAxi_wa_ready = _T ? 1'h0 : _GEN_408; // @[Conditional.scala 40:58 axi.scala 101:18]
  assign io_flashAxi_wd_ready = _T ? 1'h0 : _GEN_407; // @[Conditional.scala 40:58 axi.scala 102:18]
  assign io_flashAxi_wr_valid = _T ? 1'h0 : _GEN_406; // @[Conditional.scala 40:58 axi.scala 103:18]
  assign io_flashAxi_wr_bits_id = _T ? 4'h0 : _GEN_405; // @[Conditional.scala 40:58 axi.scala 58:23]
  assign io_flashAxi_wr_bits_resp = _T ? 2'h0 : _GEN_404; // @[Conditional.scala 40:58 axi.scala 58:23]
  assign io_flashAxi_ra_ready = _T ? 1'h0 : _GEN_403; // @[Conditional.scala 40:58 axi.scala 104:18]
  assign io_flashAxi_rd_valid = _T ? 1'h0 : _GEN_402; // @[Conditional.scala 40:58 axi.scala 105:18]
  assign io_flashAxi_rd_bits_id = _T ? 4'h0 : _GEN_401; // @[Conditional.scala 40:58 axi.scala 68:23]
  assign io_flashAxi_rd_bits_data = _T ? 64'h0 : _GEN_400; // @[Conditional.scala 40:58 axi.scala 68:23]
  assign io_flashAxi_rd_bits_resp = _T ? 2'h0 : _GEN_399; // @[Conditional.scala 40:58 axi.scala 68:23]
  assign io_flashAxi_rd_bits_last = _T ? 1'h0 : _GEN_398; // @[Conditional.scala 40:58 axi.scala 68:23]
  assign io_memAxi_wa_ready = _T ? 1'h0 : _GEN_386; // @[Conditional.scala 40:58 axi.scala 101:18]
  assign io_memAxi_wd_ready = _T ? 1'h0 : _GEN_379; // @[Conditional.scala 40:58 axi.scala 102:18]
  assign io_memAxi_ra_ready = _T ? 1'h0 : _GEN_370; // @[Conditional.scala 40:58 axi.scala 104:18]
  assign io_memAxi_rd_valid = _T ? 1'h0 : _GEN_362; // @[Conditional.scala 40:58 axi.scala 105:18]
  assign io_memAxi_rd_bits_data = _T ? 64'h0 : _GEN_360; // @[Conditional.scala 40:58 axi.scala 68:23]
  assign io_memAxi_rd_bits_last = _T ? 1'h0 : _GEN_358; // @[Conditional.scala 40:58 axi.scala 68:23]
  assign io_mmioAxi_wa_ready = _T ? 1'h0 : _GEN_419; // @[Conditional.scala 40:58 axi.scala 101:18]
  assign io_mmioAxi_wd_ready = _T ? 1'h0 : _GEN_418; // @[Conditional.scala 40:58 axi.scala 102:18]
  assign io_mmioAxi_wr_valid = _T ? 1'h0 : _GEN_417; // @[Conditional.scala 40:58 axi.scala 103:18]
  assign io_mmioAxi_wr_bits_id = _T ? 4'h0 : _GEN_416; // @[Conditional.scala 40:58 axi.scala 58:23]
  assign io_mmioAxi_wr_bits_resp = _T ? 2'h0 : _GEN_415; // @[Conditional.scala 40:58 axi.scala 58:23]
  assign io_mmioAxi_ra_ready = _T ? 1'h0 : _GEN_414; // @[Conditional.scala 40:58 axi.scala 104:18]
  assign io_mmioAxi_rd_valid = _T ? 1'h0 : _GEN_413; // @[Conditional.scala 40:58 axi.scala 105:18]
  assign io_mmioAxi_rd_bits_id = _T ? 4'h0 : _GEN_412; // @[Conditional.scala 40:58 axi.scala 68:23]
  assign io_mmioAxi_rd_bits_data = _T ? 64'h0 : _GEN_411; // @[Conditional.scala 40:58 axi.scala 68:23]
  assign io_mmioAxi_rd_bits_resp = _T ? 2'h0 : _GEN_410; // @[Conditional.scala 40:58 axi.scala 68:23]
  assign io_mmioAxi_rd_bits_last = _T ? 1'h0 : _GEN_409; // @[Conditional.scala 40:58 axi.scala 68:23]
  assign io_outAxi_wa_valid = _T ? 1'h0 : _GEN_385; // @[Conditional.scala 40:58 axi.scala 83:18]
  assign io_outAxi_wa_bits_id = _T ? 4'h0 : _GEN_384; // @[Conditional.scala 40:58 axi.scala 41:23]
  assign io_outAxi_wa_bits_addr = _T ? 32'h0 : _GEN_383; // @[Conditional.scala 40:58 axi.scala 41:23]
  assign io_outAxi_wa_bits_len = _T ? 8'h0 : _GEN_382; // @[Conditional.scala 40:58 axi.scala 41:23]
  assign io_outAxi_wa_bits_size = _T ? 3'h0 : _GEN_381; // @[Conditional.scala 40:58 axi.scala 41:23]
  assign io_outAxi_wa_bits_burst = _T ? 2'h0 : _GEN_380; // @[Conditional.scala 40:58 axi.scala 41:23]
  assign io_outAxi_wd_valid = _T ? 1'h0 : _GEN_378; // @[Conditional.scala 40:58 axi.scala 84:18]
  assign io_outAxi_wd_bits_data = _T ? 64'h0 : _GEN_377; // @[Conditional.scala 40:58 axi.scala 50:23]
  assign io_outAxi_wd_bits_strb = _T ? 8'h0 : _GEN_376; // @[Conditional.scala 40:58 axi.scala 50:23]
  assign io_outAxi_wd_bits_last = _T ? 1'h0 : _GEN_375; // @[Conditional.scala 40:58 axi.scala 50:23]
  assign io_outAxi_wr_ready = _T | _GEN_374; // @[Conditional.scala 40:58 crossbar.scala 29:24]
  assign io_outAxi_ra_valid = _T ? 1'h0 : _GEN_369; // @[Conditional.scala 40:58 axi.scala 86:18]
  assign io_outAxi_ra_bits_id = _T ? 4'h0 : _GEN_368; // @[Conditional.scala 40:58 axi.scala 41:23]
  assign io_outAxi_ra_bits_addr = _T ? 32'h0 : _GEN_367; // @[Conditional.scala 40:58 axi.scala 41:23]
  assign io_outAxi_ra_bits_len = _T ? 8'h0 : _GEN_366; // @[Conditional.scala 40:58 axi.scala 41:23]
  assign io_outAxi_ra_bits_size = _T ? 3'h0 : _GEN_365; // @[Conditional.scala 40:58 axi.scala 41:23]
  assign io_outAxi_ra_bits_burst = _T ? 2'h0 : _GEN_364; // @[Conditional.scala 40:58 axi.scala 41:23]
  assign io_outAxi_rd_ready = _T ? 1'h0 : _GEN_363; // @[Conditional.scala 40:58 axi.scala 87:18]
  always @(posedge clock) begin
    if (reset) begin // @[crossbar.scala 20:24]
      state <= 4'h0; // @[crossbar.scala 20:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_selectMem) begin // @[crossbar.scala 42:31]
        state <= 4'h1; // @[crossbar.scala 43:23]
      end else if (io_memAxi_ra_valid | io_memAxi_wa_valid) begin // @[crossbar.scala 45:65]
        state <= 4'h1; // @[crossbar.scala 46:23]
      end else begin
        state <= _GEN_2;
      end
    end else if (_T_3) begin // @[Conditional.scala 39:67]
      if (selectMem_r & ~io_selectMem) begin // @[crossbar.scala 56:47]
        state <= 4'h0; // @[crossbar.scala 57:23]
      end else begin
        state <= _GEN_6;
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      state <= _GEN_38;
    end else begin
      state <= _GEN_269;
    end
    if (reset) begin // @[crossbar.scala 22:30]
      selectMem_r <= 1'h0; // @[crossbar.scala 22:30]
    end else if (_T) begin // @[Conditional.scala 40:58]
      selectMem_r <= _GEN_5;
    end else if (_T_3) begin // @[Conditional.scala 39:67]
      if (selectMem_r & ~io_selectMem) begin // @[crossbar.scala 56:47]
        selectMem_r <= 1'h0; // @[crossbar.scala 58:29]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      selectMem_r <= _GEN_39;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  selectMem_r = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_FetchCrossBar(
  input         clock,
  input         reset,
  input  [31:0] io_instIO_addr,
  output [63:0] io_instIO_inst,
  input         io_instIO_arvalid,
  output        io_instIO_rvalid,
  output [31:0] io_icRead_addr,
  input  [63:0] io_icRead_inst,
  output        io_icRead_arvalid,
  input         io_icRead_rvalid,
  output [31:0] io_flashRead_addr,
  input  [63:0] io_flashRead_rdata,
  input         io_flashRead_rvalid,
  output [4:0]  io_flashRead_dc_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  pre_mem; // @[fetch.scala 18:26]
  wire  inp_mem = io_instIO_addr[31]; // @[fetch.scala 19:33]
  wire [4:0] _GEN_2 = inp_mem ? 5'h0 : 5'h7; // @[fetch.scala 28:22 fetch.scala 22:26 fetch.scala 32:34]
  assign io_instIO_inst = pre_mem ? io_icRead_inst : io_flashRead_rdata; // @[fetch.scala 38:18 fetch.scala 39:25 fetch.scala 42:25]
  assign io_instIO_rvalid = pre_mem ? io_icRead_rvalid : io_flashRead_rvalid; // @[fetch.scala 38:18 fetch.scala 40:26 fetch.scala 43:26]
  assign io_icRead_addr = io_instIO_addr; // @[fetch.scala 23:25]
  assign io_icRead_arvalid = io_instIO_arvalid & inp_mem; // @[fetch.scala 26:28 fetch.scala 24:25]
  assign io_flashRead_addr = io_instIO_addr; // @[fetch.scala 20:25]
  assign io_flashRead_dc_mode = io_instIO_arvalid ? _GEN_2 : 5'h0; // @[fetch.scala 26:28 fetch.scala 22:26]
  always @(posedge clock) begin
    if (reset) begin // @[fetch.scala 18:26]
      pre_mem <= 1'h0; // @[fetch.scala 18:26]
    end else if (io_instIO_arvalid) begin // @[fetch.scala 26:28]
      pre_mem <= inp_mem; // @[fetch.scala 27:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pre_mem = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_Splite64to32(
  input         clock,
  input         reset,
  input  [31:0] io_data_in_addr,
  output [63:0] io_data_in_rdata,
  output        io_data_in_rvalid,
  input  [4:0]  io_data_in_dc_mode,
  output [31:0] io_data_out_addr,
  input  [63:0] io_data_out_rdata,
  input         io_data_out_rvalid,
  output [4:0]  io_data_out_dc_mode,
  input         io_data_out_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] data_buf; // @[toaxi.scala 16:27]
  reg [31:0] addr_r; // @[toaxi.scala 18:25]
  reg  is_64; // @[toaxi.scala 19:24]
  reg  busy; // @[toaxi.scala 20:23]
  reg  state; // @[toaxi.scala 21:24]
  wire  hs_out = io_data_out_dc_mode != 5'h0 & io_data_out_ready; // @[toaxi.scala 22:53]
  wire [31:0] io_data_in_rdata_hi = io_data_out_rdata[31:0]; // @[toaxi.scala 25:57]
  wire [63:0] _io_data_in_rdata_T = {io_data_in_rdata_hi,data_buf}; // @[Cat.scala 30:58]
  wire  _T = ~state; // @[Conditional.scala 37:30]
  wire [28:0] io_data_out_addr_hi = io_data_in_addr[31:3]; // @[toaxi.scala 30:60]
  wire [31:0] _io_data_out_addr_T = {io_data_out_addr_hi,3'h0}; // @[Cat.scala 30:58]
  wire  _GEN_0 = hs_out ? 1'h0 : is_64; // @[toaxi.scala 37:39 toaxi.scala 38:31 toaxi.scala 19:24]
  wire  _GEN_1 = hs_out & io_data_out_dc_mode != 5'h7 | state; // @[toaxi.scala 33:68 toaxi.scala 34:31 toaxi.scala 21:24]
  wire  _GEN_3 = hs_out & io_data_out_dc_mode != 5'h7 | _GEN_0; // @[toaxi.scala 33:68 toaxi.scala 36:31]
  wire  _GEN_4 = io_data_in_rvalid ? 1'h0 : busy; // @[toaxi.scala 40:46 toaxi.scala 41:26 toaxi.scala 20:23]
  wire  _GEN_5 = io_data_in_dc_mode != 5'h0 | _GEN_4; // @[toaxi.scala 28:54 toaxi.scala 29:26]
  wire [31:0] _GEN_6 = io_data_in_dc_mode != 5'h0 ? _io_data_out_addr_T : 32'h0; // @[toaxi.scala 28:54 toaxi.scala 30:38 toaxi.scala 23:108]
  wire [4:0] _GEN_7 = io_data_in_dc_mode != 5'h0 ? 5'h16 : 5'h0; // @[toaxi.scala 28:54 toaxi.scala 31:41 toaxi.scala 23:77]
  wire  _GEN_12 = busy & io_data_out_rvalid; // @[toaxi.scala 43:27 toaxi.scala 44:39 toaxi.scala 24:52]
  wire [63:0] _GEN_13 = io_data_out_rvalid ? io_data_out_rdata : {{32'd0}, data_buf}; // @[toaxi.scala 48:37 toaxi.scala 49:26 toaxi.scala 16:27]
  wire [31:0] _io_data_out_addr_T_2 = addr_r + 32'h4; // @[toaxi.scala 51:40]
  wire [63:0] _GEN_15 = state ? _GEN_13 : {{32'd0}, data_buf}; // @[Conditional.scala 39:67 toaxi.scala 16:27]
  wire [31:0] _GEN_16 = state ? _io_data_out_addr_T_2 : 32'h0; // @[Conditional.scala 39:67 toaxi.scala 51:30 toaxi.scala 23:108]
  wire [4:0] _GEN_17 = state ? 5'h16 : 5'h0; // @[Conditional.scala 39:67 toaxi.scala 52:33 toaxi.scala 23:77]
  wire [63:0] _GEN_27 = _T ? {{32'd0}, data_buf} : _GEN_15; // @[Conditional.scala 40:58 toaxi.scala 16:27]
  assign io_data_in_rdata = is_64 ? _io_data_in_rdata_T : io_data_out_rdata; // @[toaxi.scala 25:28]
  assign io_data_in_rvalid = _T & _GEN_12; // @[Conditional.scala 40:58 toaxi.scala 24:52]
  assign io_data_out_addr = _T ? _GEN_6 : _GEN_16; // @[Conditional.scala 40:58]
  assign io_data_out_dc_mode = _T ? _GEN_7 : _GEN_17; // @[Conditional.scala 40:58]
  always @(posedge clock) begin
    if (reset) begin // @[toaxi.scala 16:27]
      data_buf <= 32'h0; // @[toaxi.scala 16:27]
    end else begin
      data_buf <= _GEN_27[31:0];
    end
    if (reset) begin // @[toaxi.scala 18:25]
      addr_r <= 32'h0; // @[toaxi.scala 18:25]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_data_in_dc_mode != 5'h0) begin // @[toaxi.scala 28:54]
        if (hs_out & io_data_out_dc_mode != 5'h7) begin // @[toaxi.scala 33:68]
          addr_r <= _io_data_out_addr_T; // @[toaxi.scala 35:32]
        end
      end
    end
    if (reset) begin // @[toaxi.scala 19:24]
      is_64 <= 1'h0; // @[toaxi.scala 19:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_data_in_dc_mode != 5'h0) begin // @[toaxi.scala 28:54]
        is_64 <= _GEN_3;
      end
    end
    if (reset) begin // @[toaxi.scala 20:23]
      busy <= 1'h0; // @[toaxi.scala 20:23]
    end else if (_T) begin // @[Conditional.scala 40:58]
      busy <= _GEN_5;
    end
    if (reset) begin // @[toaxi.scala 21:24]
      state <= 1'h0; // @[toaxi.scala 21:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_data_in_dc_mode != 5'h0) begin // @[toaxi.scala 28:54]
        state <= _GEN_1;
      end
    end else if (state) begin // @[Conditional.scala 39:67]
      if (hs_out) begin // @[toaxi.scala 53:25]
        state <= 1'h0; // @[toaxi.scala 54:23]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_buf = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  addr_r = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  is_64 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_MemCrossBar(
  input         clock,
  input         reset,
  input  [31:0] io_dataRW_addr,
  output [63:0] io_dataRW_rdata,
  output        io_dataRW_rvalid,
  input  [63:0] io_dataRW_wdata,
  input  [4:0]  io_dataRW_dc_mode,
  input  [4:0]  io_dataRW_amo,
  output        io_dataRW_ready,
  output [31:0] io_mmio_addr,
  input  [63:0] io_mmio_rdata,
  input         io_mmio_rvalid,
  output [63:0] io_mmio_wdata,
  output [4:0]  io_mmio_dc_mode,
  input         io_mmio_ready,
  output [31:0] io_dcRW_addr,
  input  [63:0] io_dcRW_rdata,
  input         io_dcRW_rvalid,
  output [63:0] io_dcRW_wdata,
  output [4:0]  io_dcRW_dc_mode,
  output [4:0]  io_dcRW_amo,
  input         io_dcRW_ready,
  output [31:0] io_clintIO_addr,
  input  [63:0] io_clintIO_rdata,
  output [63:0] io_clintIO_wdata,
  output        io_clintIO_wvalid,
  output [31:0] io_plicIO_addr,
  input  [63:0] io_plicIO_rdata,
  output [63:0] io_plicIO_wdata,
  output        io_plicIO_wvalid,
  output        io_plicIO_arvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] pre_type; // @[memory.scala 23:30]
  reg [63:0] data_r; // @[memory.scala 24:30]
  reg  data_valid; // @[memory.scala 25:30]
  wire  is_clint = io_dataRW_addr == 32'h200bff8 | io_dataRW_addr == 32'h2004000 | io_dataRW_addr == 32'h2000000; // @[memory.scala 27:79]
  wire  is_plic = io_dataRW_addr >= 32'hc000000 & io_dataRW_addr <= 32'hfffffff; // @[memory.scala 28:51]
  wire  inp_mem = io_dataRW_addr[31]; // @[memory.scala 29:37]
  wire [4:0] _GEN_1 = inp_mem ? io_dataRW_dc_mode : 5'h0; // @[memory.scala 58:28 memory.scala 60:29 memory.scala 37:21]
  wire  _GEN_2 = inp_mem ? io_dcRW_ready : io_mmio_ready; // @[memory.scala 58:28 memory.scala 61:29 memory.scala 65:29]
  wire [4:0] _GEN_3 = inp_mem ? 5'h0 : io_dataRW_dc_mode; // @[memory.scala 58:28 memory.scala 38:21 memory.scala 64:29]
  wire  _GEN_5 = is_plic & io_dataRW_dc_mode[2]; // @[memory.scala 52:28 memory.scala 54:33 memory.scala 45:23]
  wire  _GEN_6 = is_plic & io_dataRW_dc_mode[3]; // @[memory.scala 52:28 memory.scala 55:33 memory.scala 44:23]
  wire  _GEN_8 = is_plic | data_valid; // @[memory.scala 52:28 memory.scala 57:33 memory.scala 25:30]
  wire [4:0] _GEN_9 = is_plic ? 5'h0 : _GEN_1; // @[memory.scala 52:28 memory.scala 37:21]
  wire  _GEN_10 = is_plic ? 1'h0 : _GEN_2; // @[memory.scala 52:28 memory.scala 42:21]
  wire [4:0] _GEN_11 = is_plic ? 5'h0 : _GEN_3; // @[memory.scala 52:28 memory.scala 38:21]
  wire  _GEN_13 = is_clint & io_dataRW_dc_mode[3]; // @[memory.scala 47:23 memory.scala 49:33 memory.scala 43:23]
  wire  _GEN_15 = is_clint | _GEN_8; // @[memory.scala 47:23 memory.scala 51:33]
  wire  _GEN_16 = is_clint ? 1'h0 : _GEN_5; // @[memory.scala 47:23 memory.scala 45:23]
  wire  _GEN_17 = is_clint ? 1'h0 : _GEN_6; // @[memory.scala 47:23 memory.scala 44:23]
  wire [4:0] _GEN_18 = is_clint ? 5'h0 : _GEN_9; // @[memory.scala 47:23 memory.scala 37:21]
  wire  _GEN_19 = is_clint ? 1'h0 : _GEN_10; // @[memory.scala 47:23 memory.scala 42:21]
  wire [4:0] _GEN_20 = is_clint ? 5'h0 : _GEN_11; // @[memory.scala 47:23 memory.scala 38:21]
  wire [63:0] _GEN_30 = pre_type == 2'h0 ? io_mmio_rdata : 64'h0; // @[memory.scala 75:33 memory.scala 76:29 memory.scala 79:29]
  wire  _GEN_31 = pre_type == 2'h0 & io_mmio_rvalid; // @[memory.scala 75:33 memory.scala 77:29 memory.scala 80:29]
  wire [63:0] _GEN_32 = pre_type == 2'h1 ? io_dcRW_rdata : _GEN_30; // @[memory.scala 72:33 memory.scala 73:29]
  wire  _GEN_33 = pre_type == 2'h1 ? io_dcRW_rvalid : _GEN_31; // @[memory.scala 72:33 memory.scala 74:29]
  assign io_dataRW_rdata = (pre_type == 2'h2 | pre_type == 2'h3) & data_valid ? data_r : _GEN_32; // @[memory.scala 68:63 memory.scala 69:29]
  assign io_dataRW_rvalid = (pre_type == 2'h2 | pre_type == 2'h3) & data_valid | _GEN_33; // @[memory.scala 68:63 memory.scala 70:29]
  assign io_dataRW_ready = io_dataRW_dc_mode != 5'h0 & _GEN_19; // @[memory.scala 46:41 memory.scala 42:21]
  assign io_mmio_addr = io_dataRW_addr; // @[memory.scala 30:21]
  assign io_mmio_wdata = io_dataRW_wdata; // @[memory.scala 31:21]
  assign io_mmio_dc_mode = io_dataRW_dc_mode != 5'h0 ? _GEN_20 : 5'h0; // @[memory.scala 46:41 memory.scala 38:21]
  assign io_dcRW_addr = io_dataRW_addr; // @[memory.scala 32:21]
  assign io_dcRW_wdata = io_dataRW_wdata; // @[memory.scala 33:21]
  assign io_dcRW_dc_mode = io_dataRW_dc_mode != 5'h0 ? _GEN_18 : 5'h0; // @[memory.scala 46:41 memory.scala 37:21]
  assign io_dcRW_amo = io_dataRW_amo; // @[memory.scala 34:21]
  assign io_clintIO_addr = io_dataRW_addr; // @[memory.scala 35:24]
  assign io_clintIO_wdata = io_dataRW_wdata; // @[memory.scala 36:24]
  assign io_clintIO_wvalid = io_dataRW_dc_mode != 5'h0 & _GEN_13; // @[memory.scala 46:41 memory.scala 43:23]
  assign io_plicIO_addr = io_dataRW_addr; // @[memory.scala 40:21]
  assign io_plicIO_wdata = io_dataRW_wdata; // @[memory.scala 41:21]
  assign io_plicIO_wvalid = io_dataRW_dc_mode != 5'h0 & _GEN_17; // @[memory.scala 46:41 memory.scala 44:23]
  assign io_plicIO_arvalid = io_dataRW_dc_mode != 5'h0 & _GEN_16; // @[memory.scala 46:41 memory.scala 45:23]
  always @(posedge clock) begin
    if (reset) begin // @[memory.scala 23:30]
      pre_type <= 2'h0; // @[memory.scala 23:30]
    end else if (io_dataRW_dc_mode != 5'h0) begin // @[memory.scala 46:41]
      if (is_clint) begin // @[memory.scala 47:23]
        pre_type <= 2'h2; // @[memory.scala 48:33]
      end else if (is_plic) begin // @[memory.scala 52:28]
        pre_type <= 2'h3; // @[memory.scala 53:33]
      end else begin
        pre_type <= {{1'd0}, inp_mem};
      end
    end
    if (reset) begin // @[memory.scala 24:30]
      data_r <= 64'h0; // @[memory.scala 24:30]
    end else if (io_dataRW_dc_mode != 5'h0) begin // @[memory.scala 46:41]
      if (is_clint) begin // @[memory.scala 47:23]
        data_r <= io_clintIO_rdata; // @[memory.scala 50:33]
      end else if (is_plic) begin // @[memory.scala 52:28]
        data_r <= io_plicIO_rdata; // @[memory.scala 56:33]
      end
    end
    if (reset) begin // @[memory.scala 25:30]
      data_valid <= 1'h0; // @[memory.scala 25:30]
    end else if ((pre_type == 2'h2 | pre_type == 2'h3) & data_valid) begin // @[memory.scala 68:63]
      data_valid <= 1'h0; // @[memory.scala 71:29]
    end else if (io_dataRW_dc_mode != 5'h0) begin // @[memory.scala 46:41]
      data_valid <= _GEN_15;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pre_type = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  data_r = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  data_valid = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_MaxPeriodFibonacciLFSR_2(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 47:50]
  reg  state_1; // @[PRNG.scala 47:50]
  reg  state_2; // @[PRNG.scala 47:50]
  reg  state_3; // @[PRNG.scala 47:50]
  wire  _T = state_3 ^ state_2; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 69:10]
  assign io_out_1 = state_1; // @[PRNG.scala 69:10]
  assign io_out_2 = state_2; // @[PRNG.scala 69:10]
  assign io_out_3 = state_3; // @[PRNG.scala 69:10]
  always @(posedge clock) begin
    state_0 <= reset | _T; // @[PRNG.scala 47:50 PRNG.scala 47:50]
    if (reset) begin // @[PRNG.scala 47:50]
      state_1 <= 1'h0; // @[PRNG.scala 47:50]
    end else begin
      state_1 <= state_0;
    end
    if (reset) begin // @[PRNG.scala 47:50]
      state_2 <= 1'h0; // @[PRNG.scala 47:50]
    end else begin
      state_2 <= state_1;
    end
    if (reset) begin // @[PRNG.scala 47:50]
      state_3 <= 1'h0; // @[PRNG.scala 47:50]
    end else begin
      state_3 <= state_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_TLB(
  input         clock,
  input         reset,
  input  [63:0] io_va2pa_vaddr,
  input         io_va2pa_vvalid,
  output        io_va2pa_ready,
  output [31:0] io_va2pa_paddr,
  output        io_va2pa_pvalid,
  output [63:0] io_va2pa_tlb_excep_cause,
  output [63:0] io_va2pa_tlb_excep_tval,
  output        io_va2pa_tlb_excep_en,
  input  [1:0]  io_mmuState_priv,
  input  [63:0] io_mmuState_mstatus,
  input  [63:0] io_mmuState_satp,
  input         io_flush,
  output [31:0] io_dcacheRW_addr,
  input  [63:0] io_dcacheRW_rdata,
  input         io_dcacheRW_rvalid,
  output [63:0] io_dcacheRW_wdata,
  output [4:0]  io_dcacheRW_dc_mode,
  input         io_dcacheRW_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
`endif // RANDOMIZE_REG_INIT
  wire  select_prng_clock; // @[PRNG.scala 82:22]
  wire  select_prng_reset; // @[PRNG.scala 82:22]
  wire  select_prng_io_out_0; // @[PRNG.scala 82:22]
  wire  select_prng_io_out_1; // @[PRNG.scala 82:22]
  wire  select_prng_io_out_2; // @[PRNG.scala 82:22]
  wire  select_prng_io_out_3; // @[PRNG.scala 82:22]
  reg [51:0] tag_0; // @[tlb.scala 39:26]
  reg [51:0] tag_1; // @[tlb.scala 39:26]
  reg [51:0] tag_2; // @[tlb.scala 39:26]
  reg [51:0] tag_3; // @[tlb.scala 39:26]
  reg [51:0] tag_4; // @[tlb.scala 39:26]
  reg [51:0] tag_5; // @[tlb.scala 39:26]
  reg [51:0] tag_6; // @[tlb.scala 39:26]
  reg [51:0] tag_7; // @[tlb.scala 39:26]
  reg [51:0] tag_8; // @[tlb.scala 39:26]
  reg [51:0] tag_9; // @[tlb.scala 39:26]
  reg [51:0] tag_10; // @[tlb.scala 39:26]
  reg [51:0] tag_11; // @[tlb.scala 39:26]
  reg [51:0] tag_12; // @[tlb.scala 39:26]
  reg [51:0] tag_13; // @[tlb.scala 39:26]
  reg [51:0] tag_14; // @[tlb.scala 39:26]
  reg [51:0] tag_15; // @[tlb.scala 39:26]
  reg [19:0] paddr_0; // @[tlb.scala 40:26]
  reg [19:0] paddr_1; // @[tlb.scala 40:26]
  reg [19:0] paddr_2; // @[tlb.scala 40:26]
  reg [19:0] paddr_3; // @[tlb.scala 40:26]
  reg [19:0] paddr_4; // @[tlb.scala 40:26]
  reg [19:0] paddr_5; // @[tlb.scala 40:26]
  reg [19:0] paddr_6; // @[tlb.scala 40:26]
  reg [19:0] paddr_7; // @[tlb.scala 40:26]
  reg [19:0] paddr_8; // @[tlb.scala 40:26]
  reg [19:0] paddr_9; // @[tlb.scala 40:26]
  reg [19:0] paddr_10; // @[tlb.scala 40:26]
  reg [19:0] paddr_11; // @[tlb.scala 40:26]
  reg [19:0] paddr_12; // @[tlb.scala 40:26]
  reg [19:0] paddr_13; // @[tlb.scala 40:26]
  reg [19:0] paddr_14; // @[tlb.scala 40:26]
  reg [19:0] paddr_15; // @[tlb.scala 40:26]
  reg [9:0] info_0; // @[tlb.scala 41:26]
  reg [9:0] info_1; // @[tlb.scala 41:26]
  reg [9:0] info_2; // @[tlb.scala 41:26]
  reg [9:0] info_3; // @[tlb.scala 41:26]
  reg [9:0] info_4; // @[tlb.scala 41:26]
  reg [9:0] info_5; // @[tlb.scala 41:26]
  reg [9:0] info_6; // @[tlb.scala 41:26]
  reg [9:0] info_7; // @[tlb.scala 41:26]
  reg [9:0] info_8; // @[tlb.scala 41:26]
  reg [9:0] info_9; // @[tlb.scala 41:26]
  reg [9:0] info_10; // @[tlb.scala 41:26]
  reg [9:0] info_11; // @[tlb.scala 41:26]
  reg [9:0] info_12; // @[tlb.scala 41:26]
  reg [9:0] info_13; // @[tlb.scala 41:26]
  reg [9:0] info_14; // @[tlb.scala 41:26]
  reg [9:0] info_15; // @[tlb.scala 41:26]
  reg [31:0] pte_addr_0; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_1; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_2; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_3; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_4; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_5; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_6; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_7; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_8; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_9; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_10; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_11; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_12; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_13; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_14; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_15; // @[tlb.scala 42:30]
  reg [1:0] pte_level_0; // @[tlb.scala 43:30]
  reg [1:0] pte_level_1; // @[tlb.scala 43:30]
  reg [1:0] pte_level_2; // @[tlb.scala 43:30]
  reg [1:0] pte_level_3; // @[tlb.scala 43:30]
  reg [1:0] pte_level_4; // @[tlb.scala 43:30]
  reg [1:0] pte_level_5; // @[tlb.scala 43:30]
  reg [1:0] pte_level_6; // @[tlb.scala 43:30]
  reg [1:0] pte_level_7; // @[tlb.scala 43:30]
  reg [1:0] pte_level_8; // @[tlb.scala 43:30]
  reg [1:0] pte_level_9; // @[tlb.scala 43:30]
  reg [1:0] pte_level_10; // @[tlb.scala 43:30]
  reg [1:0] pte_level_11; // @[tlb.scala 43:30]
  reg [1:0] pte_level_12; // @[tlb.scala 43:30]
  reg [1:0] pte_level_13; // @[tlb.scala 43:30]
  reg [1:0] pte_level_14; // @[tlb.scala 43:30]
  reg [1:0] pte_level_15; // @[tlb.scala 43:30]
  reg  valid_0; // @[tlb.scala 44:26]
  reg  valid_1; // @[tlb.scala 44:26]
  reg  valid_2; // @[tlb.scala 44:26]
  reg  valid_3; // @[tlb.scala 44:26]
  reg  valid_4; // @[tlb.scala 44:26]
  reg  valid_5; // @[tlb.scala 44:26]
  reg  valid_6; // @[tlb.scala 44:26]
  reg  valid_7; // @[tlb.scala 44:26]
  reg  valid_8; // @[tlb.scala 44:26]
  reg  valid_9; // @[tlb.scala 44:26]
  reg  valid_10; // @[tlb.scala 44:26]
  reg  valid_11; // @[tlb.scala 44:26]
  reg  valid_12; // @[tlb.scala 44:26]
  reg  valid_13; // @[tlb.scala 44:26]
  reg  valid_14; // @[tlb.scala 44:26]
  reg  valid_15; // @[tlb.scala 44:26]
  reg [63:0] pre_addr; // @[tlb.scala 46:30]
  reg [31:0] pte_addr_r; // @[tlb.scala 47:30]
  reg [63:0] wpte_data_r; // @[tlb.scala 48:30]
  reg [4:0] dc_mode_r; // @[tlb.scala 49:30]
  reg  out_valid_r; // @[tlb.scala 51:30]
  reg [31:0] out_paddr_r; // @[tlb.scala 52:30]
  reg [63:0] out_excep_r_cause; // @[tlb.scala 53:30]
  reg [63:0] out_excep_r_tval; // @[tlb.scala 53:30]
  reg  out_excep_r_en; // @[tlb.scala 53:30]
  wire [51:0] inp_tag = io_va2pa_vaddr[63:12]; // @[tlb.scala 58:33]
  wire [3:0] mmuMode = io_mmuState_priv == 2'h3 ? 4'h0 : io_mmuState_satp[63:60]; // @[tlb.scala 65:22]
  wire  is_Sv39 = mmuMode == 4'h8; // @[tlb.scala 66:27]
  wire [51:0] _tlb_tag_mask_T_4 = 2'h0 == pte_level_0 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_6 = 2'h1 == pte_level_0 ? 52'hffffffffffe00 : _tlb_tag_mask_T_4; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask = 2'h2 == pte_level_0 ? 52'hffffffffc0000 : _tlb_tag_mask_T_6; // @[Mux.scala 80:57]
  wire [51:0] _T_1 = inp_tag & tlb_tag_mask; // @[tlb.scala 73:24]
  wire [19:0] _GEN_2 = _T_1 == tag_0 & valid_0 ? paddr_0 : 20'h0; // @[tlb.scala 73:64 tlb.scala 75:28 tlb.scala 68:40]
  wire [9:0] _GEN_4 = _T_1 == tag_0 & valid_0 ? info_0 : 10'h0; // @[tlb.scala 73:64 tlb.scala 77:28 tlb.scala 68:86]
  wire [31:0] _GEN_5 = _T_1 == tag_0 & valid_0 ? pte_addr_0 : 32'h0; // @[tlb.scala 73:64 tlb.scala 78:31 tlb.scala 69:23]
  wire [1:0] _GEN_7 = _T_1 == tag_0 & valid_0 ? pte_level_0 : 2'h0; // @[tlb.scala 73:64 tlb.scala 80:31 tlb.scala 69:69]
  wire [51:0] _tlb_tag_mask_T_12 = 2'h0 == pte_level_1 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_14 = 2'h1 == pte_level_1 ? 52'hffffffffffe00 : _tlb_tag_mask_T_12; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_1 = 2'h2 == pte_level_1 ? 52'hffffffffc0000 : _tlb_tag_mask_T_14; // @[Mux.scala 80:57]
  wire [51:0] _T_4 = inp_tag & tlb_tag_mask_1; // @[tlb.scala 73:24]
  wire  _T_6 = _T_4 == tag_1 & valid_1; // @[tlb.scala 73:52]
  wire [19:0] _GEN_9 = _T_4 == tag_1 & valid_1 ? paddr_1 : _GEN_2; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_11 = _T_4 == tag_1 & valid_1 ? info_1 : _GEN_4; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_12 = _T_4 == tag_1 & valid_1 ? pte_addr_1 : _GEN_5; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [1:0] _GEN_14 = _T_4 == tag_1 & valid_1 ? pte_level_1 : _GEN_7; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_20 = 2'h0 == pte_level_2 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_22 = 2'h1 == pte_level_2 ? 52'hffffffffffe00 : _tlb_tag_mask_T_20; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_2 = 2'h2 == pte_level_2 ? 52'hffffffffc0000 : _tlb_tag_mask_T_22; // @[Mux.scala 80:57]
  wire [51:0] _T_7 = inp_tag & tlb_tag_mask_2; // @[tlb.scala 73:24]
  wire [19:0] _GEN_16 = _T_7 == tag_2 & valid_2 ? paddr_2 : _GEN_9; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_18 = _T_7 == tag_2 & valid_2 ? info_2 : _GEN_11; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_19 = _T_7 == tag_2 & valid_2 ? pte_addr_2 : _GEN_12; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [1:0] _GEN_20 = _T_7 == tag_2 & valid_2 ? 2'h2 : {{1'd0}, _T_6}; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_21 = _T_7 == tag_2 & valid_2 ? pte_level_2 : _GEN_14; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_28 = 2'h0 == pte_level_3 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_30 = 2'h1 == pte_level_3 ? 52'hffffffffffe00 : _tlb_tag_mask_T_28; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_3 = 2'h2 == pte_level_3 ? 52'hffffffffc0000 : _tlb_tag_mask_T_30; // @[Mux.scala 80:57]
  wire [51:0] _T_10 = inp_tag & tlb_tag_mask_3; // @[tlb.scala 73:24]
  wire [19:0] _GEN_23 = _T_10 == tag_3 & valid_3 ? paddr_3 : _GEN_16; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_25 = _T_10 == tag_3 & valid_3 ? info_3 : _GEN_18; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_26 = _T_10 == tag_3 & valid_3 ? pte_addr_3 : _GEN_19; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [1:0] _GEN_27 = _T_10 == tag_3 & valid_3 ? 2'h3 : _GEN_20; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_28 = _T_10 == tag_3 & valid_3 ? pte_level_3 : _GEN_21; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_36 = 2'h0 == pte_level_4 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_38 = 2'h1 == pte_level_4 ? 52'hffffffffffe00 : _tlb_tag_mask_T_36; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_4 = 2'h2 == pte_level_4 ? 52'hffffffffc0000 : _tlb_tag_mask_T_38; // @[Mux.scala 80:57]
  wire [51:0] _T_13 = inp_tag & tlb_tag_mask_4; // @[tlb.scala 73:24]
  wire [19:0] _GEN_30 = _T_13 == tag_4 & valid_4 ? paddr_4 : _GEN_23; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_32 = _T_13 == tag_4 & valid_4 ? info_4 : _GEN_25; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_33 = _T_13 == tag_4 & valid_4 ? pte_addr_4 : _GEN_26; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [2:0] _GEN_34 = _T_13 == tag_4 & valid_4 ? 3'h4 : {{1'd0}, _GEN_27}; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_35 = _T_13 == tag_4 & valid_4 ? pte_level_4 : _GEN_28; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_44 = 2'h0 == pte_level_5 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_46 = 2'h1 == pte_level_5 ? 52'hffffffffffe00 : _tlb_tag_mask_T_44; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_5 = 2'h2 == pte_level_5 ? 52'hffffffffc0000 : _tlb_tag_mask_T_46; // @[Mux.scala 80:57]
  wire [51:0] _T_16 = inp_tag & tlb_tag_mask_5; // @[tlb.scala 73:24]
  wire [19:0] _GEN_37 = _T_16 == tag_5 & valid_5 ? paddr_5 : _GEN_30; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_39 = _T_16 == tag_5 & valid_5 ? info_5 : _GEN_32; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_40 = _T_16 == tag_5 & valid_5 ? pte_addr_5 : _GEN_33; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [2:0] _GEN_41 = _T_16 == tag_5 & valid_5 ? 3'h5 : _GEN_34; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_42 = _T_16 == tag_5 & valid_5 ? pte_level_5 : _GEN_35; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_52 = 2'h0 == pte_level_6 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_54 = 2'h1 == pte_level_6 ? 52'hffffffffffe00 : _tlb_tag_mask_T_52; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_6 = 2'h2 == pte_level_6 ? 52'hffffffffc0000 : _tlb_tag_mask_T_54; // @[Mux.scala 80:57]
  wire [51:0] _T_19 = inp_tag & tlb_tag_mask_6; // @[tlb.scala 73:24]
  wire [19:0] _GEN_44 = _T_19 == tag_6 & valid_6 ? paddr_6 : _GEN_37; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_46 = _T_19 == tag_6 & valid_6 ? info_6 : _GEN_39; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_47 = _T_19 == tag_6 & valid_6 ? pte_addr_6 : _GEN_40; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [2:0] _GEN_48 = _T_19 == tag_6 & valid_6 ? 3'h6 : _GEN_41; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_49 = _T_19 == tag_6 & valid_6 ? pte_level_6 : _GEN_42; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_60 = 2'h0 == pte_level_7 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_62 = 2'h1 == pte_level_7 ? 52'hffffffffffe00 : _tlb_tag_mask_T_60; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_7 = 2'h2 == pte_level_7 ? 52'hffffffffc0000 : _tlb_tag_mask_T_62; // @[Mux.scala 80:57]
  wire [51:0] _T_22 = inp_tag & tlb_tag_mask_7; // @[tlb.scala 73:24]
  wire [19:0] _GEN_51 = _T_22 == tag_7 & valid_7 ? paddr_7 : _GEN_44; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_53 = _T_22 == tag_7 & valid_7 ? info_7 : _GEN_46; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_54 = _T_22 == tag_7 & valid_7 ? pte_addr_7 : _GEN_47; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [2:0] _GEN_55 = _T_22 == tag_7 & valid_7 ? 3'h7 : _GEN_48; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_56 = _T_22 == tag_7 & valid_7 ? pte_level_7 : _GEN_49; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_68 = 2'h0 == pte_level_8 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_70 = 2'h1 == pte_level_8 ? 52'hffffffffffe00 : _tlb_tag_mask_T_68; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_8 = 2'h2 == pte_level_8 ? 52'hffffffffc0000 : _tlb_tag_mask_T_70; // @[Mux.scala 80:57]
  wire [51:0] _T_25 = inp_tag & tlb_tag_mask_8; // @[tlb.scala 73:24]
  wire [19:0] _GEN_58 = _T_25 == tag_8 & valid_8 ? paddr_8 : _GEN_51; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_60 = _T_25 == tag_8 & valid_8 ? info_8 : _GEN_53; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_61 = _T_25 == tag_8 & valid_8 ? pte_addr_8 : _GEN_54; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [3:0] _GEN_62 = _T_25 == tag_8 & valid_8 ? 4'h8 : {{1'd0}, _GEN_55}; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_63 = _T_25 == tag_8 & valid_8 ? pte_level_8 : _GEN_56; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_76 = 2'h0 == pte_level_9 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_78 = 2'h1 == pte_level_9 ? 52'hffffffffffe00 : _tlb_tag_mask_T_76; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_9 = 2'h2 == pte_level_9 ? 52'hffffffffc0000 : _tlb_tag_mask_T_78; // @[Mux.scala 80:57]
  wire [51:0] _T_28 = inp_tag & tlb_tag_mask_9; // @[tlb.scala 73:24]
  wire  _GEN_64 = _T_28 == tag_9 & valid_9 | (_T_25 == tag_8 & valid_8 | (_T_22 == tag_7 & valid_7 | (_T_19 == tag_6 &
    valid_6 | (_T_16 == tag_5 & valid_5 | (_T_13 == tag_4 & valid_4 | (_T_10 == tag_3 & valid_3 | (_T_7 == tag_2 &
    valid_2 | (_T_4 == tag_1 & valid_1 | _T_1 == tag_0 & valid_0)))))))); // @[tlb.scala 73:64 tlb.scala 74:28]
  wire [19:0] _GEN_65 = _T_28 == tag_9 & valid_9 ? paddr_9 : _GEN_58; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_67 = _T_28 == tag_9 & valid_9 ? info_9 : _GEN_60; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_68 = _T_28 == tag_9 & valid_9 ? pte_addr_9 : _GEN_61; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [3:0] _GEN_69 = _T_28 == tag_9 & valid_9 ? 4'h9 : _GEN_62; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_70 = _T_28 == tag_9 & valid_9 ? pte_level_9 : _GEN_63; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_84 = 2'h0 == pte_level_10 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_86 = 2'h1 == pte_level_10 ? 52'hffffffffffe00 : _tlb_tag_mask_T_84; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_10 = 2'h2 == pte_level_10 ? 52'hffffffffc0000 : _tlb_tag_mask_T_86; // @[Mux.scala 80:57]
  wire [51:0] _T_31 = inp_tag & tlb_tag_mask_10; // @[tlb.scala 73:24]
  wire [19:0] _GEN_72 = _T_31 == tag_10 & valid_10 ? paddr_10 : _GEN_65; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_74 = _T_31 == tag_10 & valid_10 ? info_10 : _GEN_67; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_75 = _T_31 == tag_10 & valid_10 ? pte_addr_10 : _GEN_68; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [3:0] _GEN_76 = _T_31 == tag_10 & valid_10 ? 4'ha : _GEN_69; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_77 = _T_31 == tag_10 & valid_10 ? pte_level_10 : _GEN_70; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_92 = 2'h0 == pte_level_11 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_94 = 2'h1 == pte_level_11 ? 52'hffffffffffe00 : _tlb_tag_mask_T_92; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_11 = 2'h2 == pte_level_11 ? 52'hffffffffc0000 : _tlb_tag_mask_T_94; // @[Mux.scala 80:57]
  wire [51:0] _T_34 = inp_tag & tlb_tag_mask_11; // @[tlb.scala 73:24]
  wire [19:0] _GEN_79 = _T_34 == tag_11 & valid_11 ? paddr_11 : _GEN_72; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_81 = _T_34 == tag_11 & valid_11 ? info_11 : _GEN_74; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_82 = _T_34 == tag_11 & valid_11 ? pte_addr_11 : _GEN_75; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [3:0] _GEN_83 = _T_34 == tag_11 & valid_11 ? 4'hb : _GEN_76; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_84 = _T_34 == tag_11 & valid_11 ? pte_level_11 : _GEN_77; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_100 = 2'h0 == pte_level_12 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_102 = 2'h1 == pte_level_12 ? 52'hffffffffffe00 : _tlb_tag_mask_T_100; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_12 = 2'h2 == pte_level_12 ? 52'hffffffffc0000 : _tlb_tag_mask_T_102; // @[Mux.scala 80:57]
  wire [51:0] _T_37 = inp_tag & tlb_tag_mask_12; // @[tlb.scala 73:24]
  wire [19:0] _GEN_86 = _T_37 == tag_12 & valid_12 ? paddr_12 : _GEN_79; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_88 = _T_37 == tag_12 & valid_12 ? info_12 : _GEN_81; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_89 = _T_37 == tag_12 & valid_12 ? pte_addr_12 : _GEN_82; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [3:0] _GEN_90 = _T_37 == tag_12 & valid_12 ? 4'hc : _GEN_83; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_91 = _T_37 == tag_12 & valid_12 ? pte_level_12 : _GEN_84; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_108 = 2'h0 == pte_level_13 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_110 = 2'h1 == pte_level_13 ? 52'hffffffffffe00 : _tlb_tag_mask_T_108; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_13 = 2'h2 == pte_level_13 ? 52'hffffffffc0000 : _tlb_tag_mask_T_110; // @[Mux.scala 80:57]
  wire [51:0] _T_40 = inp_tag & tlb_tag_mask_13; // @[tlb.scala 73:24]
  wire [19:0] _GEN_93 = _T_40 == tag_13 & valid_13 ? paddr_13 : _GEN_86; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_95 = _T_40 == tag_13 & valid_13 ? info_13 : _GEN_88; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_96 = _T_40 == tag_13 & valid_13 ? pte_addr_13 : _GEN_89; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [3:0] _GEN_97 = _T_40 == tag_13 & valid_13 ? 4'hd : _GEN_90; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_98 = _T_40 == tag_13 & valid_13 ? pte_level_13 : _GEN_91; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_116 = 2'h0 == pte_level_14 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_118 = 2'h1 == pte_level_14 ? 52'hffffffffffe00 : _tlb_tag_mask_T_116; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_14 = 2'h2 == pte_level_14 ? 52'hffffffffc0000 : _tlb_tag_mask_T_118; // @[Mux.scala 80:57]
  wire [51:0] _T_43 = inp_tag & tlb_tag_mask_14; // @[tlb.scala 73:24]
  wire [19:0] _GEN_100 = _T_43 == tag_14 & valid_14 ? paddr_14 : _GEN_93; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_102 = _T_43 == tag_14 & valid_14 ? info_14 : _GEN_95; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_103 = _T_43 == tag_14 & valid_14 ? pte_addr_14 : _GEN_96; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [3:0] _GEN_104 = _T_43 == tag_14 & valid_14 ? 4'he : _GEN_97; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_105 = _T_43 == tag_14 & valid_14 ? pte_level_14 : _GEN_98; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_124 = 2'h0 == pte_level_15 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_126 = 2'h1 == pte_level_15 ? 52'hffffffffffe00 : _tlb_tag_mask_T_124; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_15 = 2'h2 == pte_level_15 ? 52'hffffffffc0000 : _tlb_tag_mask_T_126; // @[Mux.scala 80:57]
  wire [51:0] _T_46 = inp_tag & tlb_tag_mask_15; // @[tlb.scala 73:24]
  wire  tlbMsg_tlbHit = _T_46 == tag_15 & valid_15 | (_T_43 == tag_14 & valid_14 | (_T_40 == tag_13 & valid_13 | (_T_37
     == tag_12 & valid_12 | (_T_34 == tag_11 & valid_11 | (_T_31 == tag_10 & valid_10 | _GEN_64))))); // @[tlb.scala 73:64 tlb.scala 74:28]
  wire [19:0] tlbMsg_tlbPa = _T_46 == tag_15 & valid_15 ? paddr_15 : _GEN_100; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] tlbMsg_tlbInfo = _T_46 == tag_15 & valid_15 ? info_15 : _GEN_102; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] tlbMsg_tlbPteAddr = _T_46 == tag_15 & valid_15 ? pte_addr_15 : _GEN_103; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [3:0] tlbMsg_tlbIdx = _T_46 == tag_15 & valid_15 ? 4'hf : _GEN_104; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] tlbMsg_tlbLevel = _T_46 == tag_15 & valid_15 ? pte_level_15 : _GEN_105; // @[tlb.scala 73:64 tlb.scala 80:31]
  reg [1:0] state; // @[tlb.scala 84:24]
  reg  flush_r; // @[tlb.scala 85:26]
  wire  _T_50 = state == 2'h0; // @[tlb.scala 87:20]
  wire  _GEN_113 = state == 2'h0 ? 1'h0 : valid_0; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_114 = state == 2'h0 ? 1'h0 : valid_1; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_115 = state == 2'h0 ? 1'h0 : valid_2; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_116 = state == 2'h0 ? 1'h0 : valid_3; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_117 = state == 2'h0 ? 1'h0 : valid_4; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_118 = state == 2'h0 ? 1'h0 : valid_5; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_119 = state == 2'h0 ? 1'h0 : valid_6; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_120 = state == 2'h0 ? 1'h0 : valid_7; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_121 = state == 2'h0 ? 1'h0 : valid_8; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_122 = state == 2'h0 ? 1'h0 : valid_9; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_123 = state == 2'h0 ? 1'h0 : valid_10; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_124 = state == 2'h0 ? 1'h0 : valid_11; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_125 = state == 2'h0 ? 1'h0 : valid_12; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_126 = state == 2'h0 ? 1'h0 : valid_13; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_127 = state == 2'h0 ? 1'h0 : valid_14; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_128 = state == 2'h0 ? 1'h0 : valid_15; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_130 = io_flush | flush_r ? _GEN_113 : valid_0; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_131 = io_flush | flush_r ? _GEN_114 : valid_1; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_132 = io_flush | flush_r ? _GEN_115 : valid_2; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_133 = io_flush | flush_r ? _GEN_116 : valid_3; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_134 = io_flush | flush_r ? _GEN_117 : valid_4; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_135 = io_flush | flush_r ? _GEN_118 : valid_5; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_136 = io_flush | flush_r ? _GEN_119 : valid_6; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_137 = io_flush | flush_r ? _GEN_120 : valid_7; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_138 = io_flush | flush_r ? _GEN_121 : valid_8; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_139 = io_flush | flush_r ? _GEN_122 : valid_9; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_140 = io_flush | flush_r ? _GEN_123 : valid_10; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_141 = io_flush | flush_r ? _GEN_124 : valid_11; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_142 = io_flush | flush_r ? _GEN_125 : valid_12; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_143 = io_flush | flush_r ? _GEN_126 : valid_13; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_144 = io_flush | flush_r ? _GEN_127 : valid_14; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_145 = io_flush | flush_r ? _GEN_128 : valid_15; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  handshake = io_va2pa_vvalid & io_va2pa_ready; // @[tlb.scala 94:37]
  reg [1:0] m_type_r; // @[tlb.scala 95:27]
  wire [1:0] cur_m_type = handshake ? 2'h1 : m_type_r; // @[tlb.scala 96:25]
  wire  _ad_T = cur_m_type == 2'h3; // @[common.scala 243:20]
  wire [9:0] ad = cur_m_type == 2'h3 ? 10'hc0 : 10'h40; // @[common.scala 243:12]
  wire  _GEN_150 = io_va2pa_pvalid | io_va2pa_tlb_excep_en ? 1'h0 : out_valid_r; // @[tlb.scala 108:51 tlb.scala 109:21 tlb.scala 51:30]
  wire  _GEN_151 = io_va2pa_pvalid | io_va2pa_tlb_excep_en ? 1'h0 : out_excep_r_en; // @[tlb.scala 108:51 tlb.scala 110:24 tlb.scala 53:30]
  wire  dc_hand = io_dcacheRW_ready & io_dcacheRW_dc_mode != 5'h0; // @[tlb.scala 122:37]
  wire [24:0] _tlb_high_legal_T_2 = io_va2pa_vaddr[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire  tlb_high_legal = _tlb_high_legal_T_2 == io_va2pa_vaddr[63:39]; // @[tlb.scala 125:55]
  wire  _tlb_access_illegal_T_11 = cur_m_type == 2'h2 & ~(tlbMsg_tlbInfo[1] | io_mmuState_mstatus[19] & tlbMsg_tlbInfo[3
    ]); // @[tlb.scala 127:60]
  wire  _tlb_access_illegal_T_12 = cur_m_type == 2'h1 & ~tlbMsg_tlbInfo[3] | _tlb_access_illegal_T_11; // @[tlb.scala 126:89]
  wire  _tlb_access_illegal_T_16 = _ad_T & ~tlbMsg_tlbInfo[2]; // @[tlb.scala 128:57]
  wire  tlb_access_illegal = _tlb_access_illegal_T_12 | _tlb_access_illegal_T_16; // @[tlb.scala 127:152]
  wire [3:0] select = {select_prng_io_out_3,select_prng_io_out_2,select_prng_io_out_1,select_prng_io_out_0}; // @[PRNG.scala 86:17]
  reg [3:0] select_r; // @[tlb.scala 130:27]
  reg [7:0] offset; // @[tlb.scala 131:26]
  reg [1:0] level; // @[tlb.scala 132:26]
  reg  wpte_hs_r; // @[tlb.scala 134:28]
  wire  _T_54 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire [51:0] _paddr_mask_T_4 = 2'h0 == tlbMsg_tlbLevel ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _paddr_mask_T_6 = 2'h1 == tlbMsg_tlbLevel ? 52'hffffffffffe00 : _paddr_mask_T_4; // @[Mux.scala 80:57]
  wire [51:0] paddr_mask_hi = 2'h2 == tlbMsg_tlbLevel ? 52'hffffffffc0000 : _paddr_mask_T_6; // @[Mux.scala 80:57]
  wire [63:0] paddr_mask = {paddr_mask_hi,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _out_paddr_r_T = {tlbMsg_tlbPa, 12'h0}; // @[tlb.scala 148:93]
  wire [63:0] _out_paddr_r_T_1 = ~paddr_mask; // @[common.scala 201:19]
  wire [63:0] _out_paddr_r_T_2 = io_va2pa_vaddr & _out_paddr_r_T_1; // @[common.scala 201:17]
  wire [63:0] _GEN_1417 = {{32'd0}, _out_paddr_r_T}; // @[common.scala 201:36]
  wire [63:0] _out_paddr_r_T_3 = _GEN_1417 & paddr_mask; // @[common.scala 201:36]
  wire [63:0] _out_paddr_r_T_4 = _out_paddr_r_T_2 | _out_paddr_r_T_3; // @[common.scala 201:26]
  wire [9:0] _T_59 = ad & tlbMsg_tlbInfo; // @[tlb.scala 149:30]
  wire [9:0] wpte_data_r_lo = tlbMsg_tlbInfo | ad; // @[tlb.scala 153:84]
  wire [63:0] _wpte_data_r_T = {34'h0,tlbMsg_tlbPa,wpte_data_r_lo}; // @[Cat.scala 30:58]
  wire [9:0] _GEN_152 = 4'h0 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_0; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_153 = 4'h1 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_1; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_154 = 4'h2 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_2; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_155 = 4'h3 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_3; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_156 = 4'h4 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_4; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_157 = 4'h5 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_5; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_158 = 4'h6 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_6; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_159 = 4'h7 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_7; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_160 = 4'h8 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_8; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_161 = 4'h9 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_9; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_162 = 4'ha == tlbMsg_tlbIdx ? wpte_data_r_lo : info_10; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_163 = 4'hb == tlbMsg_tlbIdx ? wpte_data_r_lo : info_11; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_164 = 4'hc == tlbMsg_tlbIdx ? wpte_data_r_lo : info_12; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_165 = 4'hd == tlbMsg_tlbIdx ? wpte_data_r_lo : info_13; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_166 = 4'he == tlbMsg_tlbIdx ? wpte_data_r_lo : info_14; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_167 = 4'hf == tlbMsg_tlbIdx ? wpte_data_r_lo : info_15; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [1:0] _GEN_168 = _T_59 != ad & is_Sv39 ? 2'h3 : state; // @[tlb.scala 149:66 tlb.scala 150:31 tlb.scala 84:24]
  wire  _GEN_169 = _T_59 != ad & is_Sv39 ? 1'h0 : wpte_hs_r; // @[tlb.scala 149:66 tlb.scala 151:35 tlb.scala 134:28]
  wire [31:0] _GEN_170 = _T_59 != ad & is_Sv39 ? tlbMsg_tlbPteAddr : pte_addr_r; // @[tlb.scala 149:66 tlb.scala 152:37 tlb.scala 47:30]
  wire [63:0] _GEN_171 = _T_59 != ad & is_Sv39 ? _wpte_data_r_T : wpte_data_r; // @[tlb.scala 149:66 tlb.scala 153:37 tlb.scala 48:30]
  wire [9:0] _GEN_172 = _T_59 != ad & is_Sv39 ? _GEN_152 : info_0; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_173 = _T_59 != ad & is_Sv39 ? _GEN_153 : info_1; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_174 = _T_59 != ad & is_Sv39 ? _GEN_154 : info_2; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_175 = _T_59 != ad & is_Sv39 ? _GEN_155 : info_3; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_176 = _T_59 != ad & is_Sv39 ? _GEN_156 : info_4; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_177 = _T_59 != ad & is_Sv39 ? _GEN_157 : info_5; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_178 = _T_59 != ad & is_Sv39 ? _GEN_158 : info_6; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_179 = _T_59 != ad & is_Sv39 ? _GEN_159 : info_7; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_180 = _T_59 != ad & is_Sv39 ? _GEN_160 : info_8; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_181 = _T_59 != ad & is_Sv39 ? _GEN_161 : info_9; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_182 = _T_59 != ad & is_Sv39 ? _GEN_162 : info_10; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_183 = _T_59 != ad & is_Sv39 ? _GEN_163 : info_11; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_184 = _T_59 != ad & is_Sv39 ? _GEN_164 : info_12; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_185 = _T_59 != ad & is_Sv39 ? _GEN_165 : info_13; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_186 = _T_59 != ad & is_Sv39 ? _GEN_166 : info_14; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_187 = _T_59 != ad & is_Sv39 ? _GEN_167 : info_15; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [43:0] pte_addr_r_hi_hi = io_mmuState_satp[43:0]; // @[tlb.scala 166:59]
  wire [63:0] _pte_addr_r_T = {{30'd0}, io_va2pa_vaddr[63:30]}; // @[tlb.scala 166:83]
  wire [8:0] pte_addr_r_hi_lo = _pte_addr_r_T[8:0]; // @[tlb.scala 166:91]
  wire [55:0] _pte_addr_r_T_1 = {pte_addr_r_hi_hi,pte_addr_r_hi_lo,3'h0}; // @[Cat.scala 30:58]
  wire  _GEN_188 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 | _GEN_151; // @[tlb.scala 162:81 tlb.scala 164:40]
  wire [55:0] _GEN_189 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 ? {{24'd0}, pte_addr_r} : _pte_addr_r_T_1; // @[tlb.scala 162:81 tlb.scala 47:30 tlb.scala 166:36]
  wire [4:0] _GEN_190 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 ? 5'h0 : 5'h7; // @[tlb.scala 162:81 tlb.scala 138:27 tlb.scala 167:36]
  wire [7:0] _GEN_191 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 ? offset : 8'h1e; // @[tlb.scala 162:81 tlb.scala 131:26 tlb.scala 168:33]
  wire [1:0] _GEN_192 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 ? level : 2'h3; // @[tlb.scala 162:81 tlb.scala 132:26 tlb.scala 169:33]
  wire [1:0] _GEN_194 = ~tlbMsg_tlbHit ? 2'h1 : state; // @[tlb.scala 156:43 tlb.scala 84:24]
  wire [3:0] _GEN_195 = ~tlbMsg_tlbHit ? select : select_r; // @[tlb.scala 156:43 tlb.scala 158:32 tlb.scala 130:27]
  wire [1:0] _GEN_196 = ~tlbMsg_tlbHit ? 2'h1 : m_type_r; // @[tlb.scala 156:43 tlb.scala 159:32 tlb.scala 95:27]
  wire [63:0] _GEN_197 = ~tlbMsg_tlbHit ? 64'hc : out_excep_r_cause; // @[tlb.scala 156:43 tlb.scala 160:39 tlb.scala 53:30]
  wire [63:0] _GEN_198 = ~tlbMsg_tlbHit ? io_va2pa_vaddr : out_excep_r_tval; // @[tlb.scala 156:43 tlb.scala 161:39 tlb.scala 53:30]
  wire  _GEN_199 = ~tlbMsg_tlbHit ? _GEN_188 : _GEN_151; // @[tlb.scala 156:43]
  wire [55:0] _GEN_200 = ~tlbMsg_tlbHit ? _GEN_189 : {{24'd0}, pte_addr_r}; // @[tlb.scala 156:43 tlb.scala 47:30]
  wire [4:0] _GEN_201 = ~tlbMsg_tlbHit ? _GEN_190 : 5'h0; // @[tlb.scala 156:43 tlb.scala 138:27]
  wire [7:0] _GEN_202 = ~tlbMsg_tlbHit ? _GEN_191 : offset; // @[tlb.scala 156:43 tlb.scala 131:26]
  wire [1:0] _GEN_203 = ~tlbMsg_tlbHit ? _GEN_192 : level; // @[tlb.scala 156:43 tlb.scala 132:26]
  wire  _GEN_204 = tlbMsg_tlbHit | _GEN_150; // @[tlb.scala 144:42 tlb.scala 145:33]
  wire [63:0] _GEN_205 = tlbMsg_tlbHit ? _out_paddr_r_T_4 : {{32'd0}, out_paddr_r}; // @[tlb.scala 144:42 tlb.scala 148:33 tlb.scala 52:30]
  wire [1:0] _GEN_206 = tlbMsg_tlbHit ? _GEN_168 : _GEN_194; // @[tlb.scala 144:42]
  wire  _GEN_207 = tlbMsg_tlbHit ? _GEN_169 : wpte_hs_r; // @[tlb.scala 144:42 tlb.scala 134:28]
  wire [55:0] _GEN_208 = tlbMsg_tlbHit ? {{24'd0}, _GEN_170} : _GEN_200; // @[tlb.scala 144:42]
  wire [63:0] _GEN_209 = tlbMsg_tlbHit ? _GEN_171 : wpte_data_r; // @[tlb.scala 144:42 tlb.scala 48:30]
  wire [9:0] _GEN_210 = tlbMsg_tlbHit ? _GEN_172 : info_0; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_211 = tlbMsg_tlbHit ? _GEN_173 : info_1; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_212 = tlbMsg_tlbHit ? _GEN_174 : info_2; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_213 = tlbMsg_tlbHit ? _GEN_175 : info_3; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_214 = tlbMsg_tlbHit ? _GEN_176 : info_4; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_215 = tlbMsg_tlbHit ? _GEN_177 : info_5; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_216 = tlbMsg_tlbHit ? _GEN_178 : info_6; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_217 = tlbMsg_tlbHit ? _GEN_179 : info_7; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_218 = tlbMsg_tlbHit ? _GEN_180 : info_8; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_219 = tlbMsg_tlbHit ? _GEN_181 : info_9; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_220 = tlbMsg_tlbHit ? _GEN_182 : info_10; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_221 = tlbMsg_tlbHit ? _GEN_183 : info_11; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_222 = tlbMsg_tlbHit ? _GEN_184 : info_12; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_223 = tlbMsg_tlbHit ? _GEN_185 : info_13; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_224 = tlbMsg_tlbHit ? _GEN_186 : info_14; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_225 = tlbMsg_tlbHit ? _GEN_187 : info_15; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [3:0] _GEN_226 = tlbMsg_tlbHit ? select_r : _GEN_195; // @[tlb.scala 144:42 tlb.scala 130:27]
  wire [1:0] _GEN_227 = tlbMsg_tlbHit ? m_type_r : _GEN_196; // @[tlb.scala 144:42 tlb.scala 95:27]
  wire [63:0] _GEN_228 = tlbMsg_tlbHit ? out_excep_r_cause : _GEN_197; // @[tlb.scala 144:42 tlb.scala 53:30]
  wire [63:0] _GEN_229 = tlbMsg_tlbHit ? out_excep_r_tval : _GEN_198; // @[tlb.scala 144:42 tlb.scala 53:30]
  wire  _GEN_230 = tlbMsg_tlbHit ? _GEN_151 : _GEN_199; // @[tlb.scala 144:42]
  wire [4:0] _GEN_231 = tlbMsg_tlbHit ? 5'h0 : _GEN_201; // @[tlb.scala 144:42 tlb.scala 138:27]
  wire [7:0] _GEN_232 = tlbMsg_tlbHit ? offset : _GEN_202; // @[tlb.scala 144:42 tlb.scala 131:26]
  wire [1:0] _GEN_233 = tlbMsg_tlbHit ? level : _GEN_203; // @[tlb.scala 144:42 tlb.scala 132:26]
  wire  _GEN_234 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal | _GEN_230; // @[tlb.scala 140:85 tlb.scala 141:36]
  wire [63:0] _GEN_235 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? 64'hc : _GEN_228; // @[tlb.scala 140:85 tlb.scala 142:39]
  wire [63:0] _GEN_236 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? io_va2pa_vaddr : _GEN_229; // @[tlb.scala 140:85 tlb.scala 143:39]
  wire  _GEN_237 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? _GEN_150 : _GEN_204; // @[tlb.scala 140:85]
  wire [63:0] _GEN_238 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? {{32'd0}, out_paddr_r} : _GEN_205; // @[tlb.scala 140:85 tlb.scala 52:30]
  wire [1:0] _GEN_239 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? state : _GEN_206; // @[tlb.scala 140:85 tlb.scala 84:24]
  wire  _GEN_240 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? wpte_hs_r : _GEN_207; // @[tlb.scala 140:85 tlb.scala 134:28]
  wire [55:0] _GEN_241 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? {{24'd0}, pte_addr_r} : _GEN_208; // @[tlb.scala 140:85 tlb.scala 47:30]
  wire [63:0] _GEN_242 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? wpte_data_r : _GEN_209; // @[tlb.scala 140:85 tlb.scala 48:30]
  wire [9:0] _GEN_243 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_0 : _GEN_210; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_244 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_1 : _GEN_211; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_245 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_2 : _GEN_212; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_246 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_3 : _GEN_213; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_247 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_4 : _GEN_214; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_248 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_5 : _GEN_215; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_249 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_6 : _GEN_216; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_250 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_7 : _GEN_217; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_251 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_8 : _GEN_218; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_252 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_9 : _GEN_219; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_253 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_10 : _GEN_220; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_254 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_11 : _GEN_221; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_255 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_12 : _GEN_222; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_256 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_13 : _GEN_223; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_257 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_14 : _GEN_224; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_258 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_15 : _GEN_225; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [3:0] _GEN_259 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? select_r : _GEN_226; // @[tlb.scala 140:85 tlb.scala 130:27]
  wire [1:0] _GEN_260 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? m_type_r : _GEN_227; // @[tlb.scala 140:85 tlb.scala 95:27]
  wire [4:0] _GEN_261 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? 5'h0 : _GEN_231; // @[tlb.scala 140:85 tlb.scala 138:27]
  wire [7:0] _GEN_262 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? offset : _GEN_232; // @[tlb.scala 140:85 tlb.scala 131:26]
  wire [1:0] _GEN_263 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? level : _GEN_233; // @[tlb.scala 140:85 tlb.scala 132:26]
  wire [63:0] _GEN_268 = ~handshake ? {{32'd0}, out_paddr_r} : _GEN_238; // @[tlb.scala 139:33 tlb.scala 52:30]
  wire [55:0] _GEN_271 = ~handshake ? {{24'd0}, pte_addr_r} : _GEN_241; // @[tlb.scala 139:33 tlb.scala 47:30]
  wire  _T_68 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [4:0] _dc_mode_r_T = wpte_hs_r ? 5'h0 : 5'hb; // @[tlb.scala 175:33]
  wire [4:0] _GEN_294 = io_dcacheRW_ready ? 5'h0 : _dc_mode_r_T; // @[tlb.scala 176:40 tlb.scala 177:31 tlb.scala 175:27]
  wire  _GEN_295 = io_dcacheRW_ready | wpte_hs_r; // @[tlb.scala 176:40 tlb.scala 178:31 tlb.scala 134:28]
  wire [1:0] _GEN_296 = io_dcacheRW_rvalid ? 2'h0 : state; // @[tlb.scala 180:41 tlb.scala 181:27 tlb.scala 84:24]
  wire  _T_69 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire [7:0] _offset_T_1 = offset - 8'h9; // @[tlb.scala 187:39]
  wire [1:0] _level_T_1 = level - 2'h1; // @[tlb.scala 188:38]
  wire [4:0] _GEN_297 = dc_hand ? 5'h0 : dc_mode_r; // @[tlb.scala 185:30 tlb.scala 186:31 tlb.scala 49:30]
  wire [7:0] _GEN_298 = dc_hand ? _offset_T_1 : offset; // @[tlb.scala 185:30 tlb.scala 187:29 tlb.scala 131:26]
  wire [1:0] _GEN_299 = dc_hand ? _level_T_1 : level; // @[tlb.scala 185:30 tlb.scala 188:29 tlb.scala 132:26]
  wire [63:0] _T_73 = io_dcacheRW_rdata & 64'hf; // @[tlb.scala 191:31]
  wire [63:0] _T_77 = io_dcacheRW_rdata & 64'hd0; // @[tlb.scala 192:35]
  wire [43:0] pte_addr_r_hi_hi_1 = io_dcacheRW_rdata[53:10]; // @[tlb.scala 196:50]
  wire [63:0] _pte_addr_r_T_2 = pre_addr >> offset; // @[tlb.scala 196:69]
  wire [8:0] pte_addr_r_hi_lo_1 = _pte_addr_r_T_2[8:0]; // @[tlb.scala 196:79]
  wire [55:0] _pte_addr_r_T_3 = {pte_addr_r_hi_hi_1,pte_addr_r_hi_lo_1,3'h0}; // @[Cat.scala 30:58]
  wire [1:0] _GEN_300 = _T_77 != 64'h0 ? 2'h0 : state; // @[tlb.scala 192:70 tlb.scala 193:35 tlb.scala 84:24]
  wire  _GEN_301 = _T_77 != 64'h0 | _GEN_151; // @[tlb.scala 192:70 tlb.scala 194:44]
  wire [55:0] _GEN_302 = _T_77 != 64'h0 ? {{24'd0}, pte_addr_r} : _pte_addr_r_T_3; // @[tlb.scala 192:70 tlb.scala 47:30 tlb.scala 196:40]
  wire [4:0] _GEN_303 = _T_77 != 64'h0 ? _GEN_297 : 5'h7; // @[tlb.scala 192:70 tlb.scala 197:40]
  wire  _T_83 = out_excep_r_cause == 64'hc; // @[tlb.scala 199:133]
  wire  _T_87 = io_dcacheRW_rdata[4] ? io_mmuState_priv == 2'h1 & (~io_mmuState_mstatus[18] | out_excep_r_cause == 64'hc
    ) : io_mmuState_priv == 2'h0; // @[tlb.scala 199:35]
  wire  _T_106 = out_excep_r_cause == 64'hd & ~(io_dcacheRW_rdata[1] | io_mmuState_mstatus[19] & io_dcacheRW_rdata[3]); // @[tlb.scala 208:82]
  wire  _T_107 = _T_83 & ~io_dcacheRW_rdata[3] | _T_106; // @[tlb.scala 207:102]
  wire  _T_111 = out_excep_r_cause == 64'hf & ~io_dcacheRW_rdata[2]; // @[tlb.scala 209:79]
  wire  _T_112 = _T_107 | _T_111; // @[tlb.scala 208:152]
  wire [51:0] _ppn_mask_T_4 = 2'h0 == level ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _ppn_mask_T_6 = 2'h1 == level ? 52'hffffffffffe00 : _ppn_mask_T_4; // @[Mux.scala 80:57]
  wire [51:0] ppn_mask = 2'h2 == level ? 52'hffffffffc0000 : _ppn_mask_T_6; // @[Mux.scala 80:57]
  wire [51:0] _tag_T_1 = pre_addr[63:12] & ppn_mask; // @[tlb.scala 220:78]
  wire [51:0] _GEN_304 = 4'h0 == select_r ? _tag_T_1 : tag_0; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_305 = 4'h1 == select_r ? _tag_T_1 : tag_1; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_306 = 4'h2 == select_r ? _tag_T_1 : tag_2; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_307 = 4'h3 == select_r ? _tag_T_1 : tag_3; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_308 = 4'h4 == select_r ? _tag_T_1 : tag_4; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_309 = 4'h5 == select_r ? _tag_T_1 : tag_5; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_310 = 4'h6 == select_r ? _tag_T_1 : tag_6; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_311 = 4'h7 == select_r ? _tag_T_1 : tag_7; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_312 = 4'h8 == select_r ? _tag_T_1 : tag_8; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_313 = 4'h9 == select_r ? _tag_T_1 : tag_9; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_314 = 4'ha == select_r ? _tag_T_1 : tag_10; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_315 = 4'hb == select_r ? _tag_T_1 : tag_11; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_316 = 4'hc == select_r ? _tag_T_1 : tag_12; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_317 = 4'hd == select_r ? _tag_T_1 : tag_13; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_318 = 4'he == select_r ? _tag_T_1 : tag_14; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_319 = 4'hf == select_r ? _tag_T_1 : tag_15; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire  _GEN_320 = 4'h0 == select_r | _GEN_130; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_321 = 4'h1 == select_r | _GEN_131; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_322 = 4'h2 == select_r | _GEN_132; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_323 = 4'h3 == select_r | _GEN_133; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_324 = 4'h4 == select_r | _GEN_134; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_325 = 4'h5 == select_r | _GEN_135; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_326 = 4'h6 == select_r | _GEN_136; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_327 = 4'h7 == select_r | _GEN_137; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_328 = 4'h8 == select_r | _GEN_138; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_329 = 4'h9 == select_r | _GEN_139; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_330 = 4'ha == select_r | _GEN_140; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_331 = 4'hb == select_r | _GEN_141; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_332 = 4'hc == select_r | _GEN_142; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_333 = 4'hd == select_r | _GEN_143; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_334 = 4'he == select_r | _GEN_144; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_335 = 4'hf == select_r | _GEN_145; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire [51:0] _GEN_1435 = {{32'd0}, io_dcacheRW_rdata[29:10]}; // @[tlb.scala 222:53]
  wire [51:0] update_pa = _GEN_1435 & ppn_mask; // @[tlb.scala 222:53]
  wire [19:0] _GEN_336 = 4'h0 == select_r ? update_pa[19:0] : paddr_0; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_337 = 4'h1 == select_r ? update_pa[19:0] : paddr_1; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_338 = 4'h2 == select_r ? update_pa[19:0] : paddr_2; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_339 = 4'h3 == select_r ? update_pa[19:0] : paddr_3; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_340 = 4'h4 == select_r ? update_pa[19:0] : paddr_4; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_341 = 4'h5 == select_r ? update_pa[19:0] : paddr_5; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_342 = 4'h6 == select_r ? update_pa[19:0] : paddr_6; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_343 = 4'h7 == select_r ? update_pa[19:0] : paddr_7; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_344 = 4'h8 == select_r ? update_pa[19:0] : paddr_8; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_345 = 4'h9 == select_r ? update_pa[19:0] : paddr_9; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_346 = 4'ha == select_r ? update_pa[19:0] : paddr_10; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_347 = 4'hb == select_r ? update_pa[19:0] : paddr_11; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_348 = 4'hc == select_r ? update_pa[19:0] : paddr_12; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_349 = 4'hd == select_r ? update_pa[19:0] : paddr_13; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_350 = 4'he == select_r ? update_pa[19:0] : paddr_14; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_351 = 4'hf == select_r ? update_pa[19:0] : paddr_15; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [31:0] _GEN_352 = 4'h0 == select_r ? pte_addr_r : pte_addr_0; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_353 = 4'h1 == select_r ? pte_addr_r : pte_addr_1; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_354 = 4'h2 == select_r ? pte_addr_r : pte_addr_2; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_355 = 4'h3 == select_r ? pte_addr_r : pte_addr_3; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_356 = 4'h4 == select_r ? pte_addr_r : pte_addr_4; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_357 = 4'h5 == select_r ? pte_addr_r : pte_addr_5; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_358 = 4'h6 == select_r ? pte_addr_r : pte_addr_6; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_359 = 4'h7 == select_r ? pte_addr_r : pte_addr_7; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_360 = 4'h8 == select_r ? pte_addr_r : pte_addr_8; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_361 = 4'h9 == select_r ? pte_addr_r : pte_addr_9; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_362 = 4'ha == select_r ? pte_addr_r : pte_addr_10; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_363 = 4'hb == select_r ? pte_addr_r : pte_addr_11; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_364 = 4'hc == select_r ? pte_addr_r : pte_addr_12; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_365 = 4'hd == select_r ? pte_addr_r : pte_addr_13; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_366 = 4'he == select_r ? pte_addr_r : pte_addr_14; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_367 = 4'hf == select_r ? pte_addr_r : pte_addr_15; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [1:0] _GEN_368 = 4'h0 == select_r ? level : pte_level_0; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_369 = 4'h1 == select_r ? level : pte_level_1; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_370 = 4'h2 == select_r ? level : pte_level_2; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_371 = 4'h3 == select_r ? level : pte_level_3; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_372 = 4'h4 == select_r ? level : pte_level_4; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_373 = 4'h5 == select_r ? level : pte_level_5; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_374 = 4'h6 == select_r ? level : pte_level_6; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_375 = 4'h7 == select_r ? level : pte_level_7; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_376 = 4'h8 == select_r ? level : pte_level_8; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_377 = 4'h9 == select_r ? level : pte_level_9; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_378 = 4'ha == select_r ? level : pte_level_10; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_379 = 4'hb == select_r ? level : pte_level_11; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_380 = 4'hc == select_r ? level : pte_level_12; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_381 = 4'hd == select_r ? level : pte_level_13; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_382 = 4'he == select_r ? level : pte_level_14; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_383 = 4'hf == select_r ? level : pte_level_15; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [9:0] _GEN_384 = 4'h0 == select_r ? io_dcacheRW_rdata[9:0] : info_0; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_385 = 4'h1 == select_r ? io_dcacheRW_rdata[9:0] : info_1; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_386 = 4'h2 == select_r ? io_dcacheRW_rdata[9:0] : info_2; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_387 = 4'h3 == select_r ? io_dcacheRW_rdata[9:0] : info_3; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_388 = 4'h4 == select_r ? io_dcacheRW_rdata[9:0] : info_4; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_389 = 4'h5 == select_r ? io_dcacheRW_rdata[9:0] : info_5; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_390 = 4'h6 == select_r ? io_dcacheRW_rdata[9:0] : info_6; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_391 = 4'h7 == select_r ? io_dcacheRW_rdata[9:0] : info_7; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_392 = 4'h8 == select_r ? io_dcacheRW_rdata[9:0] : info_8; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_393 = 4'h9 == select_r ? io_dcacheRW_rdata[9:0] : info_9; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_394 = 4'ha == select_r ? io_dcacheRW_rdata[9:0] : info_10; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_395 = 4'hb == select_r ? io_dcacheRW_rdata[9:0] : info_11; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_396 = 4'hc == select_r ? io_dcacheRW_rdata[9:0] : info_12; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_397 = 4'hd == select_r ? io_dcacheRW_rdata[9:0] : info_13; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_398 = 4'he == select_r ? io_dcacheRW_rdata[9:0] : info_14; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_399 = 4'hf == select_r ? io_dcacheRW_rdata[9:0] : info_15; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire  _GEN_401 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     | _GEN_151; // @[tlb.scala 213:117 tlb.scala 216:40]
  wire [51:0] _GEN_402 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_0 : _GEN_304; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_403 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_1 : _GEN_305; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_404 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_2 : _GEN_306; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_405 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_3 : _GEN_307; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_406 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_4 : _GEN_308; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_407 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_5 : _GEN_309; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_408 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_6 : _GEN_310; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_409 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_7 : _GEN_311; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_410 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_8 : _GEN_312; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_411 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_9 : _GEN_313; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_412 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_10 : _GEN_314; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_413 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_11 : _GEN_315; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_414 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_12 : _GEN_316; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_415 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_13 : _GEN_317; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_416 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_14 : _GEN_318; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_417 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_15 : _GEN_319; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire  _GEN_418 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_130 : _GEN_320; // @[tlb.scala 213:117]
  wire  _GEN_419 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_131 : _GEN_321; // @[tlb.scala 213:117]
  wire  _GEN_420 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_132 : _GEN_322; // @[tlb.scala 213:117]
  wire  _GEN_421 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_133 : _GEN_323; // @[tlb.scala 213:117]
  wire  _GEN_422 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_134 : _GEN_324; // @[tlb.scala 213:117]
  wire  _GEN_423 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_135 : _GEN_325; // @[tlb.scala 213:117]
  wire  _GEN_424 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_136 : _GEN_326; // @[tlb.scala 213:117]
  wire  _GEN_425 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_137 : _GEN_327; // @[tlb.scala 213:117]
  wire  _GEN_426 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_138 : _GEN_328; // @[tlb.scala 213:117]
  wire  _GEN_427 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_139 : _GEN_329; // @[tlb.scala 213:117]
  wire  _GEN_428 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_140 : _GEN_330; // @[tlb.scala 213:117]
  wire  _GEN_429 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_141 : _GEN_331; // @[tlb.scala 213:117]
  wire  _GEN_430 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_142 : _GEN_332; // @[tlb.scala 213:117]
  wire  _GEN_431 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_143 : _GEN_333; // @[tlb.scala 213:117]
  wire  _GEN_432 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_144 : _GEN_334; // @[tlb.scala 213:117]
  wire  _GEN_433 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_145 : _GEN_335; // @[tlb.scala 213:117]
  wire [19:0] _GEN_434 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_0 : _GEN_336; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_435 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_1 : _GEN_337; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_436 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_2 : _GEN_338; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_437 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_3 : _GEN_339; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_438 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_4 : _GEN_340; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_439 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_5 : _GEN_341; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_440 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_6 : _GEN_342; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_441 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_7 : _GEN_343; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_442 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_8 : _GEN_344; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_443 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_9 : _GEN_345; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_444 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_10 : _GEN_346; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_445 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_11 : _GEN_347; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_446 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_12 : _GEN_348; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_447 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_13 : _GEN_349; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_448 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_14 : _GEN_350; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_449 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_15 : _GEN_351; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [31:0] _GEN_450 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_0 : _GEN_352; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_451 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_1 : _GEN_353; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_452 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_2 : _GEN_354; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_453 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_3 : _GEN_355; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_454 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_4 : _GEN_356; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_455 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_5 : _GEN_357; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_456 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_6 : _GEN_358; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_457 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_7 : _GEN_359; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_458 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_8 : _GEN_360; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_459 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_9 : _GEN_361; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_460 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_10 : _GEN_362; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_461 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_11 : _GEN_363; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_462 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_12 : _GEN_364; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_463 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_13 : _GEN_365; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_464 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_14 : _GEN_366; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_465 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_15 : _GEN_367; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [1:0] _GEN_466 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_0 : _GEN_368; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_467 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_1 : _GEN_369; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_468 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_2 : _GEN_370; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_469 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_3 : _GEN_371; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_470 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_4 : _GEN_372; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_471 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_5 : _GEN_373; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_472 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_6 : _GEN_374; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_473 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_7 : _GEN_375; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_474 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_8 : _GEN_376; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_475 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_9 : _GEN_377; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_476 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_10 : _GEN_378; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_477 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_11 : _GEN_379; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_478 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_12 : _GEN_380; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_479 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_13 : _GEN_381; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_480 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_14 : _GEN_382; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_481 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_15 : _GEN_383; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [9:0] _GEN_482 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_0 : _GEN_384; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_483 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_1 : _GEN_385; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_484 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_2 : _GEN_386; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_485 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_3 : _GEN_387; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_486 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_4 : _GEN_388; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_487 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_5 : _GEN_389; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_488 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_6 : _GEN_390; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_489 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_7 : _GEN_391; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_490 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_8 : _GEN_392; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_491 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_9 : _GEN_393; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_492 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_10 : _GEN_394; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_493 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_11 : _GEN_395; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_494 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_12 : _GEN_396; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_495 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_13 : _GEN_397; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_496 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_14 : _GEN_398; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_497 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_15 : _GEN_399; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire  _GEN_499 = _T_112 | _GEN_401; // @[tlb.scala 209:99 tlb.scala 212:40]
  wire [51:0] _GEN_500 = _T_112 ? tag_0 : _GEN_402; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_501 = _T_112 ? tag_1 : _GEN_403; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_502 = _T_112 ? tag_2 : _GEN_404; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_503 = _T_112 ? tag_3 : _GEN_405; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_504 = _T_112 ? tag_4 : _GEN_406; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_505 = _T_112 ? tag_5 : _GEN_407; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_506 = _T_112 ? tag_6 : _GEN_408; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_507 = _T_112 ? tag_7 : _GEN_409; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_508 = _T_112 ? tag_8 : _GEN_410; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_509 = _T_112 ? tag_9 : _GEN_411; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_510 = _T_112 ? tag_10 : _GEN_412; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_511 = _T_112 ? tag_11 : _GEN_413; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_512 = _T_112 ? tag_12 : _GEN_414; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_513 = _T_112 ? tag_13 : _GEN_415; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_514 = _T_112 ? tag_14 : _GEN_416; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_515 = _T_112 ? tag_15 : _GEN_417; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire  _GEN_516 = _T_112 ? _GEN_130 : _GEN_418; // @[tlb.scala 209:99]
  wire  _GEN_517 = _T_112 ? _GEN_131 : _GEN_419; // @[tlb.scala 209:99]
  wire  _GEN_518 = _T_112 ? _GEN_132 : _GEN_420; // @[tlb.scala 209:99]
  wire  _GEN_519 = _T_112 ? _GEN_133 : _GEN_421; // @[tlb.scala 209:99]
  wire  _GEN_520 = _T_112 ? _GEN_134 : _GEN_422; // @[tlb.scala 209:99]
  wire  _GEN_521 = _T_112 ? _GEN_135 : _GEN_423; // @[tlb.scala 209:99]
  wire  _GEN_522 = _T_112 ? _GEN_136 : _GEN_424; // @[tlb.scala 209:99]
  wire  _GEN_523 = _T_112 ? _GEN_137 : _GEN_425; // @[tlb.scala 209:99]
  wire  _GEN_524 = _T_112 ? _GEN_138 : _GEN_426; // @[tlb.scala 209:99]
  wire  _GEN_525 = _T_112 ? _GEN_139 : _GEN_427; // @[tlb.scala 209:99]
  wire  _GEN_526 = _T_112 ? _GEN_140 : _GEN_428; // @[tlb.scala 209:99]
  wire  _GEN_527 = _T_112 ? _GEN_141 : _GEN_429; // @[tlb.scala 209:99]
  wire  _GEN_528 = _T_112 ? _GEN_142 : _GEN_430; // @[tlb.scala 209:99]
  wire  _GEN_529 = _T_112 ? _GEN_143 : _GEN_431; // @[tlb.scala 209:99]
  wire  _GEN_530 = _T_112 ? _GEN_144 : _GEN_432; // @[tlb.scala 209:99]
  wire  _GEN_531 = _T_112 ? _GEN_145 : _GEN_433; // @[tlb.scala 209:99]
  wire [19:0] _GEN_532 = _T_112 ? paddr_0 : _GEN_434; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_533 = _T_112 ? paddr_1 : _GEN_435; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_534 = _T_112 ? paddr_2 : _GEN_436; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_535 = _T_112 ? paddr_3 : _GEN_437; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_536 = _T_112 ? paddr_4 : _GEN_438; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_537 = _T_112 ? paddr_5 : _GEN_439; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_538 = _T_112 ? paddr_6 : _GEN_440; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_539 = _T_112 ? paddr_7 : _GEN_441; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_540 = _T_112 ? paddr_8 : _GEN_442; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_541 = _T_112 ? paddr_9 : _GEN_443; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_542 = _T_112 ? paddr_10 : _GEN_444; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_543 = _T_112 ? paddr_11 : _GEN_445; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_544 = _T_112 ? paddr_12 : _GEN_446; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_545 = _T_112 ? paddr_13 : _GEN_447; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_546 = _T_112 ? paddr_14 : _GEN_448; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_547 = _T_112 ? paddr_15 : _GEN_449; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [31:0] _GEN_548 = _T_112 ? pte_addr_0 : _GEN_450; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_549 = _T_112 ? pte_addr_1 : _GEN_451; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_550 = _T_112 ? pte_addr_2 : _GEN_452; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_551 = _T_112 ? pte_addr_3 : _GEN_453; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_552 = _T_112 ? pte_addr_4 : _GEN_454; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_553 = _T_112 ? pte_addr_5 : _GEN_455; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_554 = _T_112 ? pte_addr_6 : _GEN_456; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_555 = _T_112 ? pte_addr_7 : _GEN_457; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_556 = _T_112 ? pte_addr_8 : _GEN_458; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_557 = _T_112 ? pte_addr_9 : _GEN_459; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_558 = _T_112 ? pte_addr_10 : _GEN_460; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_559 = _T_112 ? pte_addr_11 : _GEN_461; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_560 = _T_112 ? pte_addr_12 : _GEN_462; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_561 = _T_112 ? pte_addr_13 : _GEN_463; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_562 = _T_112 ? pte_addr_14 : _GEN_464; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_563 = _T_112 ? pte_addr_15 : _GEN_465; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [1:0] _GEN_564 = _T_112 ? pte_level_0 : _GEN_466; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_565 = _T_112 ? pte_level_1 : _GEN_467; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_566 = _T_112 ? pte_level_2 : _GEN_468; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_567 = _T_112 ? pte_level_3 : _GEN_469; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_568 = _T_112 ? pte_level_4 : _GEN_470; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_569 = _T_112 ? pte_level_5 : _GEN_471; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_570 = _T_112 ? pte_level_6 : _GEN_472; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_571 = _T_112 ? pte_level_7 : _GEN_473; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_572 = _T_112 ? pte_level_8 : _GEN_474; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_573 = _T_112 ? pte_level_9 : _GEN_475; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_574 = _T_112 ? pte_level_10 : _GEN_476; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_575 = _T_112 ? pte_level_11 : _GEN_477; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_576 = _T_112 ? pte_level_12 : _GEN_478; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_577 = _T_112 ? pte_level_13 : _GEN_479; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_578 = _T_112 ? pte_level_14 : _GEN_480; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_579 = _T_112 ? pte_level_15 : _GEN_481; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [9:0] _GEN_580 = _T_112 ? info_0 : _GEN_482; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_581 = _T_112 ? info_1 : _GEN_483; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_582 = _T_112 ? info_2 : _GEN_484; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_583 = _T_112 ? info_3 : _GEN_485; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_584 = _T_112 ? info_4 : _GEN_486; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_585 = _T_112 ? info_5 : _GEN_487; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_586 = _T_112 ? info_6 : _GEN_488; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_587 = _T_112 ? info_7 : _GEN_489; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_588 = _T_112 ? info_8 : _GEN_490; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_589 = _T_112 ? info_9 : _GEN_491; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_590 = _T_112 ? info_10 : _GEN_492; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_591 = _T_112 ? info_11 : _GEN_493; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_592 = _T_112 ? info_12 : _GEN_494; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_593 = _T_112 ? info_13 : _GEN_495; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_594 = _T_112 ? info_14 : _GEN_496; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_595 = _T_112 ? info_15 : _GEN_497; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire  _GEN_597 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] | _GEN_499; // @[tlb.scala 203:87 tlb.scala 206:40]
  wire [51:0] _GEN_598 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_0 : _GEN_500; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_599 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_1 : _GEN_501; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_600 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_2 : _GEN_502; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_601 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_3 : _GEN_503; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_602 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_4 : _GEN_504; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_603 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_5 : _GEN_505; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_604 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_6 : _GEN_506; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_605 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_7 : _GEN_507; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_606 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_8 : _GEN_508; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_607 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_9 : _GEN_509; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_608 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_10 : _GEN_510; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_609 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_11 : _GEN_511; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_610 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_12 : _GEN_512; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_611 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_13 : _GEN_513; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_612 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_14 : _GEN_514; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_613 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_15 : _GEN_515; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire  _GEN_614 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_130 : _GEN_516; // @[tlb.scala 203:87]
  wire  _GEN_615 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_131 : _GEN_517; // @[tlb.scala 203:87]
  wire  _GEN_616 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_132 : _GEN_518; // @[tlb.scala 203:87]
  wire  _GEN_617 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_133 : _GEN_519; // @[tlb.scala 203:87]
  wire  _GEN_618 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_134 : _GEN_520; // @[tlb.scala 203:87]
  wire  _GEN_619 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_135 : _GEN_521; // @[tlb.scala 203:87]
  wire  _GEN_620 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_136 : _GEN_522; // @[tlb.scala 203:87]
  wire  _GEN_621 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_137 : _GEN_523; // @[tlb.scala 203:87]
  wire  _GEN_622 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_138 : _GEN_524; // @[tlb.scala 203:87]
  wire  _GEN_623 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_139 : _GEN_525; // @[tlb.scala 203:87]
  wire  _GEN_624 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_140 : _GEN_526; // @[tlb.scala 203:87]
  wire  _GEN_625 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_141 : _GEN_527; // @[tlb.scala 203:87]
  wire  _GEN_626 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_142 : _GEN_528; // @[tlb.scala 203:87]
  wire  _GEN_627 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_143 : _GEN_529; // @[tlb.scala 203:87]
  wire  _GEN_628 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_144 : _GEN_530; // @[tlb.scala 203:87]
  wire  _GEN_629 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_145 : _GEN_531; // @[tlb.scala 203:87]
  wire [19:0] _GEN_630 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_0 : _GEN_532; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_631 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_1 : _GEN_533; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_632 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_2 : _GEN_534; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_633 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_3 : _GEN_535; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_634 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_4 : _GEN_536; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_635 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_5 : _GEN_537; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_636 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_6 : _GEN_538; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_637 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_7 : _GEN_539; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_638 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_8 : _GEN_540; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_639 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_9 : _GEN_541; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_640 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_10 : _GEN_542; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_641 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_11 : _GEN_543; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_642 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_12 : _GEN_544; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_643 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_13 : _GEN_545; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_644 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_14 : _GEN_546; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_645 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_15 : _GEN_547; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [31:0] _GEN_646 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_0 : _GEN_548; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_647 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_1 : _GEN_549; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_648 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_2 : _GEN_550; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_649 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_3 : _GEN_551; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_650 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_4 : _GEN_552; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_651 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_5 : _GEN_553; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_652 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_6 : _GEN_554; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_653 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_7 : _GEN_555; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_654 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_8 : _GEN_556; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_655 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_9 : _GEN_557; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_656 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_10 : _GEN_558; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_657 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_11 : _GEN_559; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_658 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_12 : _GEN_560; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_659 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_13 : _GEN_561; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_660 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_14 : _GEN_562; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_661 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_15 : _GEN_563; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [1:0] _GEN_662 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_0 : _GEN_564; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_663 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_1 : _GEN_565; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_664 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_2 : _GEN_566; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_665 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_3 : _GEN_567; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_666 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_4 : _GEN_568; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_667 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_5 : _GEN_569; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_668 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_6 : _GEN_570; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_669 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_7 : _GEN_571; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_670 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_8 : _GEN_572; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_671 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_9 : _GEN_573; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_672 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_10 : _GEN_574; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_673 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_11 : _GEN_575; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_674 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_12 : _GEN_576; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_675 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_13 : _GEN_577; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_676 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_14 : _GEN_578; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_677 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_15 : _GEN_579; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [9:0] _GEN_678 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_0 : _GEN_580; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_679 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_1 : _GEN_581; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_680 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_2 : _GEN_582; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_681 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_3 : _GEN_583; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_682 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_4 : _GEN_584; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_683 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_5 : _GEN_585; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_684 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_6 : _GEN_586; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_685 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_7 : _GEN_587; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_686 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_8 : _GEN_588; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_687 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_9 : _GEN_589; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_688 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_10 : _GEN_590; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_689 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_11 : _GEN_591; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_690 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_12 : _GEN_592; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_691 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_13 : _GEN_593; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_692 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_14 : _GEN_594; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_693 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_15 : _GEN_595; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire  _GEN_695 = _T_87 | _GEN_597; // @[tlb.scala 199:193 tlb.scala 202:40]
  wire [51:0] _GEN_696 = _T_87 ? tag_0 : _GEN_598; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_697 = _T_87 ? tag_1 : _GEN_599; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_698 = _T_87 ? tag_2 : _GEN_600; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_699 = _T_87 ? tag_3 : _GEN_601; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_700 = _T_87 ? tag_4 : _GEN_602; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_701 = _T_87 ? tag_5 : _GEN_603; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_702 = _T_87 ? tag_6 : _GEN_604; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_703 = _T_87 ? tag_7 : _GEN_605; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_704 = _T_87 ? tag_8 : _GEN_606; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_705 = _T_87 ? tag_9 : _GEN_607; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_706 = _T_87 ? tag_10 : _GEN_608; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_707 = _T_87 ? tag_11 : _GEN_609; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_708 = _T_87 ? tag_12 : _GEN_610; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_709 = _T_87 ? tag_13 : _GEN_611; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_710 = _T_87 ? tag_14 : _GEN_612; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_711 = _T_87 ? tag_15 : _GEN_613; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire  _GEN_712 = _T_87 ? _GEN_130 : _GEN_614; // @[tlb.scala 199:193]
  wire  _GEN_713 = _T_87 ? _GEN_131 : _GEN_615; // @[tlb.scala 199:193]
  wire  _GEN_714 = _T_87 ? _GEN_132 : _GEN_616; // @[tlb.scala 199:193]
  wire  _GEN_715 = _T_87 ? _GEN_133 : _GEN_617; // @[tlb.scala 199:193]
  wire  _GEN_716 = _T_87 ? _GEN_134 : _GEN_618; // @[tlb.scala 199:193]
  wire  _GEN_717 = _T_87 ? _GEN_135 : _GEN_619; // @[tlb.scala 199:193]
  wire  _GEN_718 = _T_87 ? _GEN_136 : _GEN_620; // @[tlb.scala 199:193]
  wire  _GEN_719 = _T_87 ? _GEN_137 : _GEN_621; // @[tlb.scala 199:193]
  wire  _GEN_720 = _T_87 ? _GEN_138 : _GEN_622; // @[tlb.scala 199:193]
  wire  _GEN_721 = _T_87 ? _GEN_139 : _GEN_623; // @[tlb.scala 199:193]
  wire  _GEN_722 = _T_87 ? _GEN_140 : _GEN_624; // @[tlb.scala 199:193]
  wire  _GEN_723 = _T_87 ? _GEN_141 : _GEN_625; // @[tlb.scala 199:193]
  wire  _GEN_724 = _T_87 ? _GEN_142 : _GEN_626; // @[tlb.scala 199:193]
  wire  _GEN_725 = _T_87 ? _GEN_143 : _GEN_627; // @[tlb.scala 199:193]
  wire  _GEN_726 = _T_87 ? _GEN_144 : _GEN_628; // @[tlb.scala 199:193]
  wire  _GEN_727 = _T_87 ? _GEN_145 : _GEN_629; // @[tlb.scala 199:193]
  wire [19:0] _GEN_728 = _T_87 ? paddr_0 : _GEN_630; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_729 = _T_87 ? paddr_1 : _GEN_631; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_730 = _T_87 ? paddr_2 : _GEN_632; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_731 = _T_87 ? paddr_3 : _GEN_633; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_732 = _T_87 ? paddr_4 : _GEN_634; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_733 = _T_87 ? paddr_5 : _GEN_635; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_734 = _T_87 ? paddr_6 : _GEN_636; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_735 = _T_87 ? paddr_7 : _GEN_637; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_736 = _T_87 ? paddr_8 : _GEN_638; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_737 = _T_87 ? paddr_9 : _GEN_639; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_738 = _T_87 ? paddr_10 : _GEN_640; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_739 = _T_87 ? paddr_11 : _GEN_641; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_740 = _T_87 ? paddr_12 : _GEN_642; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_741 = _T_87 ? paddr_13 : _GEN_643; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_742 = _T_87 ? paddr_14 : _GEN_644; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_743 = _T_87 ? paddr_15 : _GEN_645; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [31:0] _GEN_744 = _T_87 ? pte_addr_0 : _GEN_646; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_745 = _T_87 ? pte_addr_1 : _GEN_647; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_746 = _T_87 ? pte_addr_2 : _GEN_648; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_747 = _T_87 ? pte_addr_3 : _GEN_649; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_748 = _T_87 ? pte_addr_4 : _GEN_650; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_749 = _T_87 ? pte_addr_5 : _GEN_651; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_750 = _T_87 ? pte_addr_6 : _GEN_652; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_751 = _T_87 ? pte_addr_7 : _GEN_653; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_752 = _T_87 ? pte_addr_8 : _GEN_654; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_753 = _T_87 ? pte_addr_9 : _GEN_655; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_754 = _T_87 ? pte_addr_10 : _GEN_656; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_755 = _T_87 ? pte_addr_11 : _GEN_657; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_756 = _T_87 ? pte_addr_12 : _GEN_658; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_757 = _T_87 ? pte_addr_13 : _GEN_659; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_758 = _T_87 ? pte_addr_14 : _GEN_660; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_759 = _T_87 ? pte_addr_15 : _GEN_661; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [1:0] _GEN_760 = _T_87 ? pte_level_0 : _GEN_662; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_761 = _T_87 ? pte_level_1 : _GEN_663; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_762 = _T_87 ? pte_level_2 : _GEN_664; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_763 = _T_87 ? pte_level_3 : _GEN_665; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_764 = _T_87 ? pte_level_4 : _GEN_666; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_765 = _T_87 ? pte_level_5 : _GEN_667; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_766 = _T_87 ? pte_level_6 : _GEN_668; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_767 = _T_87 ? pte_level_7 : _GEN_669; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_768 = _T_87 ? pte_level_8 : _GEN_670; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_769 = _T_87 ? pte_level_9 : _GEN_671; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_770 = _T_87 ? pte_level_10 : _GEN_672; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_771 = _T_87 ? pte_level_11 : _GEN_673; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_772 = _T_87 ? pte_level_12 : _GEN_674; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_773 = _T_87 ? pte_level_13 : _GEN_675; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_774 = _T_87 ? pte_level_14 : _GEN_676; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_775 = _T_87 ? pte_level_15 : _GEN_677; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [9:0] _GEN_776 = _T_87 ? info_0 : _GEN_678; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_777 = _T_87 ? info_1 : _GEN_679; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_778 = _T_87 ? info_2 : _GEN_680; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_779 = _T_87 ? info_3 : _GEN_681; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_780 = _T_87 ? info_4 : _GEN_682; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_781 = _T_87 ? info_5 : _GEN_683; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_782 = _T_87 ? info_6 : _GEN_684; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_783 = _T_87 ? info_7 : _GEN_685; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_784 = _T_87 ? info_8 : _GEN_686; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_785 = _T_87 ? info_9 : _GEN_687; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_786 = _T_87 ? info_10 : _GEN_688; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_787 = _T_87 ? info_11 : _GEN_689; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_788 = _T_87 ? info_12 : _GEN_690; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_789 = _T_87 ? info_13 : _GEN_691; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_790 = _T_87 ? info_14 : _GEN_692; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_791 = _T_87 ? info_15 : _GEN_693; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [1:0] _GEN_792 = _T_73 == 64'h1 ? _GEN_300 : 2'h0; // @[tlb.scala 191:76]
  wire  _GEN_793 = _T_73 == 64'h1 ? _GEN_301 : _GEN_695; // @[tlb.scala 191:76]
  wire [55:0] _GEN_794 = _T_73 == 64'h1 ? _GEN_302 : {{24'd0}, pte_addr_r}; // @[tlb.scala 191:76 tlb.scala 47:30]
  wire [4:0] _GEN_795 = _T_73 == 64'h1 ? _GEN_303 : _GEN_297; // @[tlb.scala 191:76]
  wire [51:0] _GEN_796 = _T_73 == 64'h1 ? tag_0 : _GEN_696; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_797 = _T_73 == 64'h1 ? tag_1 : _GEN_697; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_798 = _T_73 == 64'h1 ? tag_2 : _GEN_698; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_799 = _T_73 == 64'h1 ? tag_3 : _GEN_699; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_800 = _T_73 == 64'h1 ? tag_4 : _GEN_700; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_801 = _T_73 == 64'h1 ? tag_5 : _GEN_701; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_802 = _T_73 == 64'h1 ? tag_6 : _GEN_702; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_803 = _T_73 == 64'h1 ? tag_7 : _GEN_703; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_804 = _T_73 == 64'h1 ? tag_8 : _GEN_704; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_805 = _T_73 == 64'h1 ? tag_9 : _GEN_705; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_806 = _T_73 == 64'h1 ? tag_10 : _GEN_706; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_807 = _T_73 == 64'h1 ? tag_11 : _GEN_707; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_808 = _T_73 == 64'h1 ? tag_12 : _GEN_708; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_809 = _T_73 == 64'h1 ? tag_13 : _GEN_709; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_810 = _T_73 == 64'h1 ? tag_14 : _GEN_710; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_811 = _T_73 == 64'h1 ? tag_15 : _GEN_711; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire  _GEN_812 = _T_73 == 64'h1 ? _GEN_130 : _GEN_712; // @[tlb.scala 191:76]
  wire  _GEN_813 = _T_73 == 64'h1 ? _GEN_131 : _GEN_713; // @[tlb.scala 191:76]
  wire  _GEN_814 = _T_73 == 64'h1 ? _GEN_132 : _GEN_714; // @[tlb.scala 191:76]
  wire  _GEN_815 = _T_73 == 64'h1 ? _GEN_133 : _GEN_715; // @[tlb.scala 191:76]
  wire  _GEN_816 = _T_73 == 64'h1 ? _GEN_134 : _GEN_716; // @[tlb.scala 191:76]
  wire  _GEN_817 = _T_73 == 64'h1 ? _GEN_135 : _GEN_717; // @[tlb.scala 191:76]
  wire  _GEN_818 = _T_73 == 64'h1 ? _GEN_136 : _GEN_718; // @[tlb.scala 191:76]
  wire  _GEN_819 = _T_73 == 64'h1 ? _GEN_137 : _GEN_719; // @[tlb.scala 191:76]
  wire  _GEN_820 = _T_73 == 64'h1 ? _GEN_138 : _GEN_720; // @[tlb.scala 191:76]
  wire  _GEN_821 = _T_73 == 64'h1 ? _GEN_139 : _GEN_721; // @[tlb.scala 191:76]
  wire  _GEN_822 = _T_73 == 64'h1 ? _GEN_140 : _GEN_722; // @[tlb.scala 191:76]
  wire  _GEN_823 = _T_73 == 64'h1 ? _GEN_141 : _GEN_723; // @[tlb.scala 191:76]
  wire  _GEN_824 = _T_73 == 64'h1 ? _GEN_142 : _GEN_724; // @[tlb.scala 191:76]
  wire  _GEN_825 = _T_73 == 64'h1 ? _GEN_143 : _GEN_725; // @[tlb.scala 191:76]
  wire  _GEN_826 = _T_73 == 64'h1 ? _GEN_144 : _GEN_726; // @[tlb.scala 191:76]
  wire  _GEN_827 = _T_73 == 64'h1 ? _GEN_145 : _GEN_727; // @[tlb.scala 191:76]
  wire [19:0] _GEN_828 = _T_73 == 64'h1 ? paddr_0 : _GEN_728; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_829 = _T_73 == 64'h1 ? paddr_1 : _GEN_729; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_830 = _T_73 == 64'h1 ? paddr_2 : _GEN_730; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_831 = _T_73 == 64'h1 ? paddr_3 : _GEN_731; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_832 = _T_73 == 64'h1 ? paddr_4 : _GEN_732; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_833 = _T_73 == 64'h1 ? paddr_5 : _GEN_733; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_834 = _T_73 == 64'h1 ? paddr_6 : _GEN_734; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_835 = _T_73 == 64'h1 ? paddr_7 : _GEN_735; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_836 = _T_73 == 64'h1 ? paddr_8 : _GEN_736; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_837 = _T_73 == 64'h1 ? paddr_9 : _GEN_737; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_838 = _T_73 == 64'h1 ? paddr_10 : _GEN_738; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_839 = _T_73 == 64'h1 ? paddr_11 : _GEN_739; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_840 = _T_73 == 64'h1 ? paddr_12 : _GEN_740; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_841 = _T_73 == 64'h1 ? paddr_13 : _GEN_741; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_842 = _T_73 == 64'h1 ? paddr_14 : _GEN_742; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_843 = _T_73 == 64'h1 ? paddr_15 : _GEN_743; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [31:0] _GEN_844 = _T_73 == 64'h1 ? pte_addr_0 : _GEN_744; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_845 = _T_73 == 64'h1 ? pte_addr_1 : _GEN_745; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_846 = _T_73 == 64'h1 ? pte_addr_2 : _GEN_746; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_847 = _T_73 == 64'h1 ? pte_addr_3 : _GEN_747; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_848 = _T_73 == 64'h1 ? pte_addr_4 : _GEN_748; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_849 = _T_73 == 64'h1 ? pte_addr_5 : _GEN_749; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_850 = _T_73 == 64'h1 ? pte_addr_6 : _GEN_750; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_851 = _T_73 == 64'h1 ? pte_addr_7 : _GEN_751; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_852 = _T_73 == 64'h1 ? pte_addr_8 : _GEN_752; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_853 = _T_73 == 64'h1 ? pte_addr_9 : _GEN_753; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_854 = _T_73 == 64'h1 ? pte_addr_10 : _GEN_754; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_855 = _T_73 == 64'h1 ? pte_addr_11 : _GEN_755; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_856 = _T_73 == 64'h1 ? pte_addr_12 : _GEN_756; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_857 = _T_73 == 64'h1 ? pte_addr_13 : _GEN_757; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_858 = _T_73 == 64'h1 ? pte_addr_14 : _GEN_758; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_859 = _T_73 == 64'h1 ? pte_addr_15 : _GEN_759; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [1:0] _GEN_860 = _T_73 == 64'h1 ? pte_level_0 : _GEN_760; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_861 = _T_73 == 64'h1 ? pte_level_1 : _GEN_761; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_862 = _T_73 == 64'h1 ? pte_level_2 : _GEN_762; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_863 = _T_73 == 64'h1 ? pte_level_3 : _GEN_763; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_864 = _T_73 == 64'h1 ? pte_level_4 : _GEN_764; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_865 = _T_73 == 64'h1 ? pte_level_5 : _GEN_765; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_866 = _T_73 == 64'h1 ? pte_level_6 : _GEN_766; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_867 = _T_73 == 64'h1 ? pte_level_7 : _GEN_767; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_868 = _T_73 == 64'h1 ? pte_level_8 : _GEN_768; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_869 = _T_73 == 64'h1 ? pte_level_9 : _GEN_769; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_870 = _T_73 == 64'h1 ? pte_level_10 : _GEN_770; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_871 = _T_73 == 64'h1 ? pte_level_11 : _GEN_771; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_872 = _T_73 == 64'h1 ? pte_level_12 : _GEN_772; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_873 = _T_73 == 64'h1 ? pte_level_13 : _GEN_773; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_874 = _T_73 == 64'h1 ? pte_level_14 : _GEN_774; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_875 = _T_73 == 64'h1 ? pte_level_15 : _GEN_775; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [9:0] _GEN_876 = _T_73 == 64'h1 ? info_0 : _GEN_776; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_877 = _T_73 == 64'h1 ? info_1 : _GEN_777; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_878 = _T_73 == 64'h1 ? info_2 : _GEN_778; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_879 = _T_73 == 64'h1 ? info_3 : _GEN_779; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_880 = _T_73 == 64'h1 ? info_4 : _GEN_780; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_881 = _T_73 == 64'h1 ? info_5 : _GEN_781; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_882 = _T_73 == 64'h1 ? info_6 : _GEN_782; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_883 = _T_73 == 64'h1 ? info_7 : _GEN_783; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_884 = _T_73 == 64'h1 ? info_8 : _GEN_784; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_885 = _T_73 == 64'h1 ? info_9 : _GEN_785; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_886 = _T_73 == 64'h1 ? info_10 : _GEN_786; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_887 = _T_73 == 64'h1 ? info_11 : _GEN_787; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_888 = _T_73 == 64'h1 ? info_12 : _GEN_788; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_889 = _T_73 == 64'h1 ? info_13 : _GEN_789; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_890 = _T_73 == 64'h1 ? info_14 : _GEN_790; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_891 = _T_73 == 64'h1 ? info_15 : _GEN_791; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [1:0] _GEN_892 = io_dcacheRW_rvalid ? _GEN_792 : state; // @[tlb.scala 190:41 tlb.scala 84:24]
  wire  _GEN_893 = io_dcacheRW_rvalid ? _GEN_793 : _GEN_151; // @[tlb.scala 190:41]
  wire [55:0] _GEN_894 = io_dcacheRW_rvalid ? _GEN_794 : {{24'd0}, pte_addr_r}; // @[tlb.scala 190:41 tlb.scala 47:30]
  wire [4:0] _GEN_895 = io_dcacheRW_rvalid ? _GEN_795 : _GEN_297; // @[tlb.scala 190:41]
  wire [51:0] _GEN_896 = io_dcacheRW_rvalid ? _GEN_796 : tag_0; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_897 = io_dcacheRW_rvalid ? _GEN_797 : tag_1; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_898 = io_dcacheRW_rvalid ? _GEN_798 : tag_2; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_899 = io_dcacheRW_rvalid ? _GEN_799 : tag_3; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_900 = io_dcacheRW_rvalid ? _GEN_800 : tag_4; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_901 = io_dcacheRW_rvalid ? _GEN_801 : tag_5; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_902 = io_dcacheRW_rvalid ? _GEN_802 : tag_6; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_903 = io_dcacheRW_rvalid ? _GEN_803 : tag_7; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_904 = io_dcacheRW_rvalid ? _GEN_804 : tag_8; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_905 = io_dcacheRW_rvalid ? _GEN_805 : tag_9; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_906 = io_dcacheRW_rvalid ? _GEN_806 : tag_10; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_907 = io_dcacheRW_rvalid ? _GEN_807 : tag_11; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_908 = io_dcacheRW_rvalid ? _GEN_808 : tag_12; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_909 = io_dcacheRW_rvalid ? _GEN_809 : tag_13; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_910 = io_dcacheRW_rvalid ? _GEN_810 : tag_14; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_911 = io_dcacheRW_rvalid ? _GEN_811 : tag_15; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire  _GEN_912 = io_dcacheRW_rvalid ? _GEN_812 : _GEN_130; // @[tlb.scala 190:41]
  wire  _GEN_913 = io_dcacheRW_rvalid ? _GEN_813 : _GEN_131; // @[tlb.scala 190:41]
  wire  _GEN_914 = io_dcacheRW_rvalid ? _GEN_814 : _GEN_132; // @[tlb.scala 190:41]
  wire  _GEN_915 = io_dcacheRW_rvalid ? _GEN_815 : _GEN_133; // @[tlb.scala 190:41]
  wire  _GEN_916 = io_dcacheRW_rvalid ? _GEN_816 : _GEN_134; // @[tlb.scala 190:41]
  wire  _GEN_917 = io_dcacheRW_rvalid ? _GEN_817 : _GEN_135; // @[tlb.scala 190:41]
  wire  _GEN_918 = io_dcacheRW_rvalid ? _GEN_818 : _GEN_136; // @[tlb.scala 190:41]
  wire  _GEN_919 = io_dcacheRW_rvalid ? _GEN_819 : _GEN_137; // @[tlb.scala 190:41]
  wire  _GEN_920 = io_dcacheRW_rvalid ? _GEN_820 : _GEN_138; // @[tlb.scala 190:41]
  wire  _GEN_921 = io_dcacheRW_rvalid ? _GEN_821 : _GEN_139; // @[tlb.scala 190:41]
  wire  _GEN_922 = io_dcacheRW_rvalid ? _GEN_822 : _GEN_140; // @[tlb.scala 190:41]
  wire  _GEN_923 = io_dcacheRW_rvalid ? _GEN_823 : _GEN_141; // @[tlb.scala 190:41]
  wire  _GEN_924 = io_dcacheRW_rvalid ? _GEN_824 : _GEN_142; // @[tlb.scala 190:41]
  wire  _GEN_925 = io_dcacheRW_rvalid ? _GEN_825 : _GEN_143; // @[tlb.scala 190:41]
  wire  _GEN_926 = io_dcacheRW_rvalid ? _GEN_826 : _GEN_144; // @[tlb.scala 190:41]
  wire  _GEN_927 = io_dcacheRW_rvalid ? _GEN_827 : _GEN_145; // @[tlb.scala 190:41]
  wire [19:0] _GEN_928 = io_dcacheRW_rvalid ? _GEN_828 : paddr_0; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_929 = io_dcacheRW_rvalid ? _GEN_829 : paddr_1; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_930 = io_dcacheRW_rvalid ? _GEN_830 : paddr_2; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_931 = io_dcacheRW_rvalid ? _GEN_831 : paddr_3; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_932 = io_dcacheRW_rvalid ? _GEN_832 : paddr_4; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_933 = io_dcacheRW_rvalid ? _GEN_833 : paddr_5; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_934 = io_dcacheRW_rvalid ? _GEN_834 : paddr_6; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_935 = io_dcacheRW_rvalid ? _GEN_835 : paddr_7; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_936 = io_dcacheRW_rvalid ? _GEN_836 : paddr_8; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_937 = io_dcacheRW_rvalid ? _GEN_837 : paddr_9; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_938 = io_dcacheRW_rvalid ? _GEN_838 : paddr_10; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_939 = io_dcacheRW_rvalid ? _GEN_839 : paddr_11; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_940 = io_dcacheRW_rvalid ? _GEN_840 : paddr_12; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_941 = io_dcacheRW_rvalid ? _GEN_841 : paddr_13; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_942 = io_dcacheRW_rvalid ? _GEN_842 : paddr_14; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_943 = io_dcacheRW_rvalid ? _GEN_843 : paddr_15; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [31:0] _GEN_944 = io_dcacheRW_rvalid ? _GEN_844 : pte_addr_0; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_945 = io_dcacheRW_rvalid ? _GEN_845 : pte_addr_1; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_946 = io_dcacheRW_rvalid ? _GEN_846 : pte_addr_2; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_947 = io_dcacheRW_rvalid ? _GEN_847 : pte_addr_3; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_948 = io_dcacheRW_rvalid ? _GEN_848 : pte_addr_4; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_949 = io_dcacheRW_rvalid ? _GEN_849 : pte_addr_5; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_950 = io_dcacheRW_rvalid ? _GEN_850 : pte_addr_6; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_951 = io_dcacheRW_rvalid ? _GEN_851 : pte_addr_7; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_952 = io_dcacheRW_rvalid ? _GEN_852 : pte_addr_8; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_953 = io_dcacheRW_rvalid ? _GEN_853 : pte_addr_9; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_954 = io_dcacheRW_rvalid ? _GEN_854 : pte_addr_10; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_955 = io_dcacheRW_rvalid ? _GEN_855 : pte_addr_11; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_956 = io_dcacheRW_rvalid ? _GEN_856 : pte_addr_12; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_957 = io_dcacheRW_rvalid ? _GEN_857 : pte_addr_13; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_958 = io_dcacheRW_rvalid ? _GEN_858 : pte_addr_14; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_959 = io_dcacheRW_rvalid ? _GEN_859 : pte_addr_15; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [1:0] _GEN_960 = io_dcacheRW_rvalid ? _GEN_860 : pte_level_0; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_961 = io_dcacheRW_rvalid ? _GEN_861 : pte_level_1; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_962 = io_dcacheRW_rvalid ? _GEN_862 : pte_level_2; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_963 = io_dcacheRW_rvalid ? _GEN_863 : pte_level_3; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_964 = io_dcacheRW_rvalid ? _GEN_864 : pte_level_4; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_965 = io_dcacheRW_rvalid ? _GEN_865 : pte_level_5; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_966 = io_dcacheRW_rvalid ? _GEN_866 : pte_level_6; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_967 = io_dcacheRW_rvalid ? _GEN_867 : pte_level_7; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_968 = io_dcacheRW_rvalid ? _GEN_868 : pte_level_8; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_969 = io_dcacheRW_rvalid ? _GEN_869 : pte_level_9; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_970 = io_dcacheRW_rvalid ? _GEN_870 : pte_level_10; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_971 = io_dcacheRW_rvalid ? _GEN_871 : pte_level_11; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_972 = io_dcacheRW_rvalid ? _GEN_872 : pte_level_12; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_973 = io_dcacheRW_rvalid ? _GEN_873 : pte_level_13; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_974 = io_dcacheRW_rvalid ? _GEN_874 : pte_level_14; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_975 = io_dcacheRW_rvalid ? _GEN_875 : pte_level_15; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [9:0] _GEN_976 = io_dcacheRW_rvalid ? _GEN_876 : info_0; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_977 = io_dcacheRW_rvalid ? _GEN_877 : info_1; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_978 = io_dcacheRW_rvalid ? _GEN_878 : info_2; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_979 = io_dcacheRW_rvalid ? _GEN_879 : info_3; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_980 = io_dcacheRW_rvalid ? _GEN_880 : info_4; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_981 = io_dcacheRW_rvalid ? _GEN_881 : info_5; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_982 = io_dcacheRW_rvalid ? _GEN_882 : info_6; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_983 = io_dcacheRW_rvalid ? _GEN_883 : info_7; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_984 = io_dcacheRW_rvalid ? _GEN_884 : info_8; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_985 = io_dcacheRW_rvalid ? _GEN_885 : info_9; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_986 = io_dcacheRW_rvalid ? _GEN_886 : info_10; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_987 = io_dcacheRW_rvalid ? _GEN_887 : info_11; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_988 = io_dcacheRW_rvalid ? _GEN_888 : info_12; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_989 = io_dcacheRW_rvalid ? _GEN_889 : info_13; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_990 = io_dcacheRW_rvalid ? _GEN_890 : info_14; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_991 = io_dcacheRW_rvalid ? _GEN_891 : info_15; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [4:0] _GEN_992 = _T_69 ? _GEN_895 : dc_mode_r; // @[Conditional.scala 39:67 tlb.scala 49:30]
  wire [7:0] _GEN_993 = _T_69 ? _GEN_298 : offset; // @[Conditional.scala 39:67 tlb.scala 131:26]
  wire [1:0] _GEN_994 = _T_69 ? _GEN_299 : level; // @[Conditional.scala 39:67 tlb.scala 132:26]
  wire [1:0] _GEN_995 = _T_69 ? _GEN_892 : state; // @[Conditional.scala 39:67 tlb.scala 84:24]
  wire  _GEN_996 = _T_69 ? _GEN_893 : _GEN_151; // @[Conditional.scala 39:67]
  wire [55:0] _GEN_997 = _T_69 ? _GEN_894 : {{24'd0}, pte_addr_r}; // @[Conditional.scala 39:67 tlb.scala 47:30]
  wire [51:0] _GEN_998 = _T_69 ? _GEN_896 : tag_0; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_999 = _T_69 ? _GEN_897 : tag_1; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1000 = _T_69 ? _GEN_898 : tag_2; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1001 = _T_69 ? _GEN_899 : tag_3; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1002 = _T_69 ? _GEN_900 : tag_4; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1003 = _T_69 ? _GEN_901 : tag_5; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1004 = _T_69 ? _GEN_902 : tag_6; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1005 = _T_69 ? _GEN_903 : tag_7; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1006 = _T_69 ? _GEN_904 : tag_8; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1007 = _T_69 ? _GEN_905 : tag_9; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1008 = _T_69 ? _GEN_906 : tag_10; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1009 = _T_69 ? _GEN_907 : tag_11; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1010 = _T_69 ? _GEN_908 : tag_12; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1011 = _T_69 ? _GEN_909 : tag_13; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1012 = _T_69 ? _GEN_910 : tag_14; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1013 = _T_69 ? _GEN_911 : tag_15; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire  _GEN_1014 = _T_69 ? _GEN_912 : _GEN_130; // @[Conditional.scala 39:67]
  wire  _GEN_1015 = _T_69 ? _GEN_913 : _GEN_131; // @[Conditional.scala 39:67]
  wire  _GEN_1016 = _T_69 ? _GEN_914 : _GEN_132; // @[Conditional.scala 39:67]
  wire  _GEN_1017 = _T_69 ? _GEN_915 : _GEN_133; // @[Conditional.scala 39:67]
  wire  _GEN_1018 = _T_69 ? _GEN_916 : _GEN_134; // @[Conditional.scala 39:67]
  wire  _GEN_1019 = _T_69 ? _GEN_917 : _GEN_135; // @[Conditional.scala 39:67]
  wire  _GEN_1020 = _T_69 ? _GEN_918 : _GEN_136; // @[Conditional.scala 39:67]
  wire  _GEN_1021 = _T_69 ? _GEN_919 : _GEN_137; // @[Conditional.scala 39:67]
  wire  _GEN_1022 = _T_69 ? _GEN_920 : _GEN_138; // @[Conditional.scala 39:67]
  wire  _GEN_1023 = _T_69 ? _GEN_921 : _GEN_139; // @[Conditional.scala 39:67]
  wire  _GEN_1024 = _T_69 ? _GEN_922 : _GEN_140; // @[Conditional.scala 39:67]
  wire  _GEN_1025 = _T_69 ? _GEN_923 : _GEN_141; // @[Conditional.scala 39:67]
  wire  _GEN_1026 = _T_69 ? _GEN_924 : _GEN_142; // @[Conditional.scala 39:67]
  wire  _GEN_1027 = _T_69 ? _GEN_925 : _GEN_143; // @[Conditional.scala 39:67]
  wire  _GEN_1028 = _T_69 ? _GEN_926 : _GEN_144; // @[Conditional.scala 39:67]
  wire  _GEN_1029 = _T_69 ? _GEN_927 : _GEN_145; // @[Conditional.scala 39:67]
  wire [19:0] _GEN_1030 = _T_69 ? _GEN_928 : paddr_0; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1031 = _T_69 ? _GEN_929 : paddr_1; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1032 = _T_69 ? _GEN_930 : paddr_2; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1033 = _T_69 ? _GEN_931 : paddr_3; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1034 = _T_69 ? _GEN_932 : paddr_4; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1035 = _T_69 ? _GEN_933 : paddr_5; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1036 = _T_69 ? _GEN_934 : paddr_6; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1037 = _T_69 ? _GEN_935 : paddr_7; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1038 = _T_69 ? _GEN_936 : paddr_8; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1039 = _T_69 ? _GEN_937 : paddr_9; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1040 = _T_69 ? _GEN_938 : paddr_10; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1041 = _T_69 ? _GEN_939 : paddr_11; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1042 = _T_69 ? _GEN_940 : paddr_12; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1043 = _T_69 ? _GEN_941 : paddr_13; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1044 = _T_69 ? _GEN_942 : paddr_14; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1045 = _T_69 ? _GEN_943 : paddr_15; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [31:0] _GEN_1046 = _T_69 ? _GEN_944 : pte_addr_0; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1047 = _T_69 ? _GEN_945 : pte_addr_1; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1048 = _T_69 ? _GEN_946 : pte_addr_2; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1049 = _T_69 ? _GEN_947 : pte_addr_3; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1050 = _T_69 ? _GEN_948 : pte_addr_4; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1051 = _T_69 ? _GEN_949 : pte_addr_5; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1052 = _T_69 ? _GEN_950 : pte_addr_6; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1053 = _T_69 ? _GEN_951 : pte_addr_7; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1054 = _T_69 ? _GEN_952 : pte_addr_8; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1055 = _T_69 ? _GEN_953 : pte_addr_9; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1056 = _T_69 ? _GEN_954 : pte_addr_10; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1057 = _T_69 ? _GEN_955 : pte_addr_11; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1058 = _T_69 ? _GEN_956 : pte_addr_12; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1059 = _T_69 ? _GEN_957 : pte_addr_13; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1060 = _T_69 ? _GEN_958 : pte_addr_14; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1061 = _T_69 ? _GEN_959 : pte_addr_15; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [1:0] _GEN_1062 = _T_69 ? _GEN_960 : pte_level_0; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1063 = _T_69 ? _GEN_961 : pte_level_1; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1064 = _T_69 ? _GEN_962 : pte_level_2; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1065 = _T_69 ? _GEN_963 : pte_level_3; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1066 = _T_69 ? _GEN_964 : pte_level_4; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1067 = _T_69 ? _GEN_965 : pte_level_5; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1068 = _T_69 ? _GEN_966 : pte_level_6; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1069 = _T_69 ? _GEN_967 : pte_level_7; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1070 = _T_69 ? _GEN_968 : pte_level_8; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1071 = _T_69 ? _GEN_969 : pte_level_9; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1072 = _T_69 ? _GEN_970 : pte_level_10; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1073 = _T_69 ? _GEN_971 : pte_level_11; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1074 = _T_69 ? _GEN_972 : pte_level_12; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1075 = _T_69 ? _GEN_973 : pte_level_13; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1076 = _T_69 ? _GEN_974 : pte_level_14; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1077 = _T_69 ? _GEN_975 : pte_level_15; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [9:0] _GEN_1078 = _T_69 ? _GEN_976 : info_0; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1079 = _T_69 ? _GEN_977 : info_1; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1080 = _T_69 ? _GEN_978 : info_2; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1081 = _T_69 ? _GEN_979 : info_3; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1082 = _T_69 ? _GEN_980 : info_4; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1083 = _T_69 ? _GEN_981 : info_5; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1084 = _T_69 ? _GEN_982 : info_6; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1085 = _T_69 ? _GEN_983 : info_7; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1086 = _T_69 ? _GEN_984 : info_8; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1087 = _T_69 ? _GEN_985 : info_9; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1088 = _T_69 ? _GEN_986 : info_10; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1089 = _T_69 ? _GEN_987 : info_11; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1090 = _T_69 ? _GEN_988 : info_12; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1091 = _T_69 ? _GEN_989 : info_13; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1092 = _T_69 ? _GEN_990 : info_14; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1093 = _T_69 ? _GEN_991 : info_15; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [55:0] _GEN_1100 = _T_68 ? {{24'd0}, pte_addr_r} : _GEN_997; // @[Conditional.scala 39:67 tlb.scala 47:30]
  wire [63:0] _GEN_1202 = _T_54 ? _GEN_268 : {{32'd0}, out_paddr_r}; // @[Conditional.scala 40:58 tlb.scala 52:30]
  wire [55:0] _GEN_1205 = _T_54 ? _GEN_271 : _GEN_1100; // @[Conditional.scala 40:58]
  wire [63:0] _GEN_1312 = is_Sv39 | state != 2'h0 ? _GEN_1202 : io_va2pa_vaddr; // @[tlb.scala 135:37 tlb.scala 233:21]
  wire [55:0] _GEN_1315 = is_Sv39 | state != 2'h0 ? _GEN_1205 : {{24'd0}, pte_addr_r}; // @[tlb.scala 135:37 tlb.scala 47:30]
  ysyx_210539_MaxPeriodFibonacciLFSR_2 select_prng ( // @[PRNG.scala 82:22]
    .clock(select_prng_clock),
    .reset(select_prng_reset),
    .io_out_0(select_prng_io_out_0),
    .io_out_1(select_prng_io_out_1),
    .io_out_2(select_prng_io_out_2),
    .io_out_3(select_prng_io_out_3)
  );
  assign io_va2pa_ready = io_va2pa_vvalid & _T_50 & ~io_flush & ~flush_r; // @[tlb.scala 98:74]
  assign io_va2pa_paddr = out_paddr_r; // @[tlb.scala 113:20]
  assign io_va2pa_pvalid = out_valid_r; // @[tlb.scala 114:21]
  assign io_va2pa_tlb_excep_cause = out_excep_r_cause; // @[tlb.scala 115:24]
  assign io_va2pa_tlb_excep_tval = out_excep_r_tval; // @[tlb.scala 115:24]
  assign io_va2pa_tlb_excep_en = out_excep_r_en; // @[tlb.scala 115:24]
  assign io_dcacheRW_addr = pte_addr_r; // @[tlb.scala 117:22]
  assign io_dcacheRW_wdata = wpte_data_r; // @[tlb.scala 118:23]
  assign io_dcacheRW_dc_mode = dc_mode_r; // @[tlb.scala 119:25]
  assign select_prng_clock = clock;
  assign select_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[tlb.scala 39:26]
      tag_0 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_0 <= _GEN_998;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_1 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_1 <= _GEN_999;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_2 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_2 <= _GEN_1000;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_3 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_3 <= _GEN_1001;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_4 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_4 <= _GEN_1002;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_5 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_5 <= _GEN_1003;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_6 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_6 <= _GEN_1004;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_7 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_7 <= _GEN_1005;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_8 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_8 <= _GEN_1006;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_9 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_9 <= _GEN_1007;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_10 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_10 <= _GEN_1008;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_11 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_11 <= _GEN_1009;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_12 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_12 <= _GEN_1010;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_13 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_13 <= _GEN_1011;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_14 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_14 <= _GEN_1012;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_15 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_15 <= _GEN_1013;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_0 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_0 <= _GEN_1030;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_1 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_1 <= _GEN_1031;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_2 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_2 <= _GEN_1032;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_3 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_3 <= _GEN_1033;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_4 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_4 <= _GEN_1034;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_5 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_5 <= _GEN_1035;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_6 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_6 <= _GEN_1036;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_7 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_7 <= _GEN_1037;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_8 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_8 <= _GEN_1038;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_9 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_9 <= _GEN_1039;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_10 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_10 <= _GEN_1040;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_11 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_11 <= _GEN_1041;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_12 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_12 <= _GEN_1042;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_13 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_13 <= _GEN_1043;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_14 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_14 <= _GEN_1044;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_15 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_15 <= _GEN_1045;
        end
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_0 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_0 <= _GEN_243;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_0 <= _GEN_1078;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_1 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_1 <= _GEN_244;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_1 <= _GEN_1079;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_2 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_2 <= _GEN_245;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_2 <= _GEN_1080;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_3 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_3 <= _GEN_246;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_3 <= _GEN_1081;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_4 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_4 <= _GEN_247;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_4 <= _GEN_1082;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_5 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_5 <= _GEN_248;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_5 <= _GEN_1083;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_6 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_6 <= _GEN_249;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_6 <= _GEN_1084;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_7 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_7 <= _GEN_250;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_7 <= _GEN_1085;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_8 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_8 <= _GEN_251;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_8 <= _GEN_1086;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_9 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_9 <= _GEN_252;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_9 <= _GEN_1087;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_10 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_10 <= _GEN_253;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_10 <= _GEN_1088;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_11 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_11 <= _GEN_254;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_11 <= _GEN_1089;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_12 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_12 <= _GEN_255;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_12 <= _GEN_1090;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_13 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_13 <= _GEN_256;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_13 <= _GEN_1091;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_14 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_14 <= _GEN_257;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_14 <= _GEN_1092;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_15 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_15 <= _GEN_258;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_15 <= _GEN_1093;
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_0 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_0 <= _GEN_1046;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_1 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_1 <= _GEN_1047;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_2 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_2 <= _GEN_1048;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_3 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_3 <= _GEN_1049;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_4 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_4 <= _GEN_1050;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_5 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_5 <= _GEN_1051;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_6 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_6 <= _GEN_1052;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_7 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_7 <= _GEN_1053;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_8 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_8 <= _GEN_1054;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_9 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_9 <= _GEN_1055;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_10 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_10 <= _GEN_1056;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_11 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_11 <= _GEN_1057;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_12 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_12 <= _GEN_1058;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_13 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_13 <= _GEN_1059;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_14 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_14 <= _GEN_1060;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_15 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_15 <= _GEN_1061;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_0 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_0 <= _GEN_1062;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_1 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_1 <= _GEN_1063;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_2 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_2 <= _GEN_1064;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_3 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_3 <= _GEN_1065;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_4 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_4 <= _GEN_1066;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_5 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_5 <= _GEN_1067;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_6 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_6 <= _GEN_1068;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_7 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_7 <= _GEN_1069;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_8 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_8 <= _GEN_1070;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_9 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_9 <= _GEN_1071;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_10 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_10 <= _GEN_1072;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_11 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_11 <= _GEN_1073;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_12 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_12 <= _GEN_1074;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_13 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_13 <= _GEN_1075;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_14 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_14 <= _GEN_1076;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_15 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_15 <= _GEN_1077;
        end
      end
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_0 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_0 <= _GEN_130;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_0 <= _GEN_130;
      end else begin
        valid_0 <= _GEN_1014;
      end
    end else begin
      valid_0 <= _GEN_130;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_1 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_1 <= _GEN_131;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_1 <= _GEN_131;
      end else begin
        valid_1 <= _GEN_1015;
      end
    end else begin
      valid_1 <= _GEN_131;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_2 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_2 <= _GEN_132;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_2 <= _GEN_132;
      end else begin
        valid_2 <= _GEN_1016;
      end
    end else begin
      valid_2 <= _GEN_132;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_3 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_3 <= _GEN_133;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_3 <= _GEN_133;
      end else begin
        valid_3 <= _GEN_1017;
      end
    end else begin
      valid_3 <= _GEN_133;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_4 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_4 <= _GEN_134;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_4 <= _GEN_134;
      end else begin
        valid_4 <= _GEN_1018;
      end
    end else begin
      valid_4 <= _GEN_134;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_5 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_5 <= _GEN_135;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_5 <= _GEN_135;
      end else begin
        valid_5 <= _GEN_1019;
      end
    end else begin
      valid_5 <= _GEN_135;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_6 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_6 <= _GEN_136;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_6 <= _GEN_136;
      end else begin
        valid_6 <= _GEN_1020;
      end
    end else begin
      valid_6 <= _GEN_136;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_7 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_7 <= _GEN_137;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_7 <= _GEN_137;
      end else begin
        valid_7 <= _GEN_1021;
      end
    end else begin
      valid_7 <= _GEN_137;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_8 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_8 <= _GEN_138;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_8 <= _GEN_138;
      end else begin
        valid_8 <= _GEN_1022;
      end
    end else begin
      valid_8 <= _GEN_138;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_9 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_9 <= _GEN_139;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_9 <= _GEN_139;
      end else begin
        valid_9 <= _GEN_1023;
      end
    end else begin
      valid_9 <= _GEN_139;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_10 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_10 <= _GEN_140;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_10 <= _GEN_140;
      end else begin
        valid_10 <= _GEN_1024;
      end
    end else begin
      valid_10 <= _GEN_140;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_11 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_11 <= _GEN_141;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_11 <= _GEN_141;
      end else begin
        valid_11 <= _GEN_1025;
      end
    end else begin
      valid_11 <= _GEN_141;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_12 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_12 <= _GEN_142;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_12 <= _GEN_142;
      end else begin
        valid_12 <= _GEN_1026;
      end
    end else begin
      valid_12 <= _GEN_142;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_13 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_13 <= _GEN_143;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_13 <= _GEN_143;
      end else begin
        valid_13 <= _GEN_1027;
      end
    end else begin
      valid_13 <= _GEN_143;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_14 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_14 <= _GEN_144;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_14 <= _GEN_144;
      end else begin
        valid_14 <= _GEN_1028;
      end
    end else begin
      valid_14 <= _GEN_144;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_15 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_15 <= _GEN_145;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_15 <= _GEN_145;
      end else begin
        valid_15 <= _GEN_1029;
      end
    end else begin
      valid_15 <= _GEN_145;
    end
    if (reset) begin // @[tlb.scala 46:30]
      pre_addr <= 64'h0; // @[tlb.scala 46:30]
    end else if (handshake) begin // @[tlb.scala 101:20]
      pre_addr <= io_va2pa_vaddr; // @[tlb.scala 103:18]
    end else if (io_va2pa_ready & io_va2pa_vvalid) begin // @[tlb.scala 54:44]
      pre_addr <= io_va2pa_vaddr; // @[tlb.scala 55:18]
    end
    if (reset) begin // @[tlb.scala 47:30]
      pte_addr_r <= 32'h0; // @[tlb.scala 47:30]
    end else begin
      pte_addr_r <= _GEN_1315[31:0];
    end
    if (reset) begin // @[tlb.scala 48:30]
      wpte_data_r <= 64'h0; // @[tlb.scala 48:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          wpte_data_r <= _GEN_242;
        end
      end
    end
    if (reset) begin // @[tlb.scala 49:30]
      dc_mode_r <= 5'h0; // @[tlb.scala 49:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (~handshake) begin // @[tlb.scala 139:33]
          dc_mode_r <= 5'h0; // @[tlb.scala 138:27]
        end else begin
          dc_mode_r <= _GEN_261;
        end
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        dc_mode_r <= _GEN_294;
      end else begin
        dc_mode_r <= _GEN_992;
      end
    end
    if (reset) begin // @[tlb.scala 51:30]
      out_valid_r <= 1'h0; // @[tlb.scala 51:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (~handshake) begin // @[tlb.scala 139:33]
          out_valid_r <= _GEN_150;
        end else begin
          out_valid_r <= _GEN_237;
        end
      end else begin
        out_valid_r <= _GEN_150;
      end
    end else begin
      out_valid_r <= io_va2pa_vvalid; // @[tlb.scala 232:21]
    end
    if (reset) begin // @[tlb.scala 52:30]
      out_paddr_r <= 32'h0; // @[tlb.scala 52:30]
    end else begin
      out_paddr_r <= _GEN_1312[31:0];
    end
    if (reset) begin // @[tlb.scala 53:30]
      out_excep_r_cause <= 64'h0; // @[tlb.scala 53:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          out_excep_r_cause <= _GEN_235;
        end
      end
    end
    if (reset) begin // @[tlb.scala 53:30]
      out_excep_r_tval <= 64'h0; // @[tlb.scala 53:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          out_excep_r_tval <= _GEN_236;
        end
      end
    end
    if (reset) begin // @[tlb.scala 53:30]
      out_excep_r_en <= 1'h0; // @[tlb.scala 53:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (~handshake) begin // @[tlb.scala 139:33]
          out_excep_r_en <= _GEN_151;
        end else begin
          out_excep_r_en <= _GEN_234;
        end
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        out_excep_r_en <= _GEN_151;
      end else begin
        out_excep_r_en <= _GEN_996;
      end
    end else begin
      out_excep_r_en <= _GEN_151;
    end
    if (reset) begin // @[tlb.scala 84:24]
      state <= 2'h0; // @[tlb.scala 84:24]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          state <= _GEN_239;
        end
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        state <= _GEN_296;
      end else begin
        state <= _GEN_995;
      end
    end
    if (reset) begin // @[tlb.scala 85:26]
      flush_r <= 1'h0; // @[tlb.scala 85:26]
    end else if (io_flush | flush_r) begin // @[tlb.scala 86:30]
      if (state == 2'h0) begin // @[tlb.scala 87:30]
        flush_r <= 1'h0; // @[tlb.scala 89:21]
      end else begin
        flush_r <= 1'h1; // @[tlb.scala 91:21]
      end
    end
    if (reset) begin // @[tlb.scala 95:27]
      m_type_r <= 2'h0; // @[tlb.scala 95:27]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          m_type_r <= _GEN_260;
        end
      end
    end
    if (reset) begin // @[tlb.scala 130:27]
      select_r <= 4'h0; // @[tlb.scala 130:27]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          select_r <= _GEN_259;
        end
      end
    end
    if (reset) begin // @[tlb.scala 131:26]
      offset <= 8'h0; // @[tlb.scala 131:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          offset <= _GEN_262;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        offset <= _GEN_993;
      end
    end
    if (reset) begin // @[tlb.scala 132:26]
      level <= 2'h0; // @[tlb.scala 132:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          level <= _GEN_263;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        level <= _GEN_994;
      end
    end
    if (reset) begin // @[tlb.scala 134:28]
      wpte_hs_r <= 1'h0; // @[tlb.scala 134:28]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          wpte_hs_r <= _GEN_240;
        end
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        wpte_hs_r <= _GEN_295;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  tag_0 = _RAND_0[51:0];
  _RAND_1 = {2{`RANDOM}};
  tag_1 = _RAND_1[51:0];
  _RAND_2 = {2{`RANDOM}};
  tag_2 = _RAND_2[51:0];
  _RAND_3 = {2{`RANDOM}};
  tag_3 = _RAND_3[51:0];
  _RAND_4 = {2{`RANDOM}};
  tag_4 = _RAND_4[51:0];
  _RAND_5 = {2{`RANDOM}};
  tag_5 = _RAND_5[51:0];
  _RAND_6 = {2{`RANDOM}};
  tag_6 = _RAND_6[51:0];
  _RAND_7 = {2{`RANDOM}};
  tag_7 = _RAND_7[51:0];
  _RAND_8 = {2{`RANDOM}};
  tag_8 = _RAND_8[51:0];
  _RAND_9 = {2{`RANDOM}};
  tag_9 = _RAND_9[51:0];
  _RAND_10 = {2{`RANDOM}};
  tag_10 = _RAND_10[51:0];
  _RAND_11 = {2{`RANDOM}};
  tag_11 = _RAND_11[51:0];
  _RAND_12 = {2{`RANDOM}};
  tag_12 = _RAND_12[51:0];
  _RAND_13 = {2{`RANDOM}};
  tag_13 = _RAND_13[51:0];
  _RAND_14 = {2{`RANDOM}};
  tag_14 = _RAND_14[51:0];
  _RAND_15 = {2{`RANDOM}};
  tag_15 = _RAND_15[51:0];
  _RAND_16 = {1{`RANDOM}};
  paddr_0 = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  paddr_1 = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  paddr_2 = _RAND_18[19:0];
  _RAND_19 = {1{`RANDOM}};
  paddr_3 = _RAND_19[19:0];
  _RAND_20 = {1{`RANDOM}};
  paddr_4 = _RAND_20[19:0];
  _RAND_21 = {1{`RANDOM}};
  paddr_5 = _RAND_21[19:0];
  _RAND_22 = {1{`RANDOM}};
  paddr_6 = _RAND_22[19:0];
  _RAND_23 = {1{`RANDOM}};
  paddr_7 = _RAND_23[19:0];
  _RAND_24 = {1{`RANDOM}};
  paddr_8 = _RAND_24[19:0];
  _RAND_25 = {1{`RANDOM}};
  paddr_9 = _RAND_25[19:0];
  _RAND_26 = {1{`RANDOM}};
  paddr_10 = _RAND_26[19:0];
  _RAND_27 = {1{`RANDOM}};
  paddr_11 = _RAND_27[19:0];
  _RAND_28 = {1{`RANDOM}};
  paddr_12 = _RAND_28[19:0];
  _RAND_29 = {1{`RANDOM}};
  paddr_13 = _RAND_29[19:0];
  _RAND_30 = {1{`RANDOM}};
  paddr_14 = _RAND_30[19:0];
  _RAND_31 = {1{`RANDOM}};
  paddr_15 = _RAND_31[19:0];
  _RAND_32 = {1{`RANDOM}};
  info_0 = _RAND_32[9:0];
  _RAND_33 = {1{`RANDOM}};
  info_1 = _RAND_33[9:0];
  _RAND_34 = {1{`RANDOM}};
  info_2 = _RAND_34[9:0];
  _RAND_35 = {1{`RANDOM}};
  info_3 = _RAND_35[9:0];
  _RAND_36 = {1{`RANDOM}};
  info_4 = _RAND_36[9:0];
  _RAND_37 = {1{`RANDOM}};
  info_5 = _RAND_37[9:0];
  _RAND_38 = {1{`RANDOM}};
  info_6 = _RAND_38[9:0];
  _RAND_39 = {1{`RANDOM}};
  info_7 = _RAND_39[9:0];
  _RAND_40 = {1{`RANDOM}};
  info_8 = _RAND_40[9:0];
  _RAND_41 = {1{`RANDOM}};
  info_9 = _RAND_41[9:0];
  _RAND_42 = {1{`RANDOM}};
  info_10 = _RAND_42[9:0];
  _RAND_43 = {1{`RANDOM}};
  info_11 = _RAND_43[9:0];
  _RAND_44 = {1{`RANDOM}};
  info_12 = _RAND_44[9:0];
  _RAND_45 = {1{`RANDOM}};
  info_13 = _RAND_45[9:0];
  _RAND_46 = {1{`RANDOM}};
  info_14 = _RAND_46[9:0];
  _RAND_47 = {1{`RANDOM}};
  info_15 = _RAND_47[9:0];
  _RAND_48 = {1{`RANDOM}};
  pte_addr_0 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  pte_addr_1 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  pte_addr_2 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  pte_addr_3 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  pte_addr_4 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  pte_addr_5 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  pte_addr_6 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  pte_addr_7 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  pte_addr_8 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  pte_addr_9 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  pte_addr_10 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  pte_addr_11 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  pte_addr_12 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  pte_addr_13 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  pte_addr_14 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  pte_addr_15 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  pte_level_0 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  pte_level_1 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  pte_level_2 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  pte_level_3 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  pte_level_4 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  pte_level_5 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  pte_level_6 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  pte_level_7 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  pte_level_8 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  pte_level_9 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  pte_level_10 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  pte_level_11 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  pte_level_12 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  pte_level_13 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  pte_level_14 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  pte_level_15 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  valid_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_4 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_5 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_6 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_7 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_8 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_9 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_10 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_11 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_12 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_13 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_14 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_15 = _RAND_95[0:0];
  _RAND_96 = {2{`RANDOM}};
  pre_addr = _RAND_96[63:0];
  _RAND_97 = {1{`RANDOM}};
  pte_addr_r = _RAND_97[31:0];
  _RAND_98 = {2{`RANDOM}};
  wpte_data_r = _RAND_98[63:0];
  _RAND_99 = {1{`RANDOM}};
  dc_mode_r = _RAND_99[4:0];
  _RAND_100 = {1{`RANDOM}};
  out_valid_r = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  out_paddr_r = _RAND_101[31:0];
  _RAND_102 = {2{`RANDOM}};
  out_excep_r_cause = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  out_excep_r_tval = _RAND_103[63:0];
  _RAND_104 = {1{`RANDOM}};
  out_excep_r_en = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  state = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  flush_r = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  m_type_r = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  select_r = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  offset = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  level = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  wpte_hs_r = _RAND_111[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_TLB_1(
  input         clock,
  input         reset,
  input  [63:0] io_va2pa_vaddr,
  input         io_va2pa_vvalid,
  input  [1:0]  io_va2pa_m_type,
  output        io_va2pa_ready,
  output [31:0] io_va2pa_paddr,
  output        io_va2pa_pvalid,
  output [63:0] io_va2pa_tlb_excep_cause,
  output [63:0] io_va2pa_tlb_excep_tval,
  output        io_va2pa_tlb_excep_en,
  input  [1:0]  io_mmuState_priv,
  input  [63:0] io_mmuState_mstatus,
  input  [63:0] io_mmuState_satp,
  input         io_flush,
  output [31:0] io_dcacheRW_addr,
  input  [63:0] io_dcacheRW_rdata,
  input         io_dcacheRW_rvalid,
  output [63:0] io_dcacheRW_wdata,
  output [4:0]  io_dcacheRW_dc_mode,
  input         io_dcacheRW_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
`endif // RANDOMIZE_REG_INIT
  wire  select_prng_clock; // @[PRNG.scala 82:22]
  wire  select_prng_reset; // @[PRNG.scala 82:22]
  wire  select_prng_io_out_0; // @[PRNG.scala 82:22]
  wire  select_prng_io_out_1; // @[PRNG.scala 82:22]
  wire  select_prng_io_out_2; // @[PRNG.scala 82:22]
  wire  select_prng_io_out_3; // @[PRNG.scala 82:22]
  reg [51:0] tag_0; // @[tlb.scala 39:26]
  reg [51:0] tag_1; // @[tlb.scala 39:26]
  reg [51:0] tag_2; // @[tlb.scala 39:26]
  reg [51:0] tag_3; // @[tlb.scala 39:26]
  reg [51:0] tag_4; // @[tlb.scala 39:26]
  reg [51:0] tag_5; // @[tlb.scala 39:26]
  reg [51:0] tag_6; // @[tlb.scala 39:26]
  reg [51:0] tag_7; // @[tlb.scala 39:26]
  reg [51:0] tag_8; // @[tlb.scala 39:26]
  reg [51:0] tag_9; // @[tlb.scala 39:26]
  reg [51:0] tag_10; // @[tlb.scala 39:26]
  reg [51:0] tag_11; // @[tlb.scala 39:26]
  reg [51:0] tag_12; // @[tlb.scala 39:26]
  reg [51:0] tag_13; // @[tlb.scala 39:26]
  reg [51:0] tag_14; // @[tlb.scala 39:26]
  reg [51:0] tag_15; // @[tlb.scala 39:26]
  reg [19:0] paddr_0; // @[tlb.scala 40:26]
  reg [19:0] paddr_1; // @[tlb.scala 40:26]
  reg [19:0] paddr_2; // @[tlb.scala 40:26]
  reg [19:0] paddr_3; // @[tlb.scala 40:26]
  reg [19:0] paddr_4; // @[tlb.scala 40:26]
  reg [19:0] paddr_5; // @[tlb.scala 40:26]
  reg [19:0] paddr_6; // @[tlb.scala 40:26]
  reg [19:0] paddr_7; // @[tlb.scala 40:26]
  reg [19:0] paddr_8; // @[tlb.scala 40:26]
  reg [19:0] paddr_9; // @[tlb.scala 40:26]
  reg [19:0] paddr_10; // @[tlb.scala 40:26]
  reg [19:0] paddr_11; // @[tlb.scala 40:26]
  reg [19:0] paddr_12; // @[tlb.scala 40:26]
  reg [19:0] paddr_13; // @[tlb.scala 40:26]
  reg [19:0] paddr_14; // @[tlb.scala 40:26]
  reg [19:0] paddr_15; // @[tlb.scala 40:26]
  reg [9:0] info_0; // @[tlb.scala 41:26]
  reg [9:0] info_1; // @[tlb.scala 41:26]
  reg [9:0] info_2; // @[tlb.scala 41:26]
  reg [9:0] info_3; // @[tlb.scala 41:26]
  reg [9:0] info_4; // @[tlb.scala 41:26]
  reg [9:0] info_5; // @[tlb.scala 41:26]
  reg [9:0] info_6; // @[tlb.scala 41:26]
  reg [9:0] info_7; // @[tlb.scala 41:26]
  reg [9:0] info_8; // @[tlb.scala 41:26]
  reg [9:0] info_9; // @[tlb.scala 41:26]
  reg [9:0] info_10; // @[tlb.scala 41:26]
  reg [9:0] info_11; // @[tlb.scala 41:26]
  reg [9:0] info_12; // @[tlb.scala 41:26]
  reg [9:0] info_13; // @[tlb.scala 41:26]
  reg [9:0] info_14; // @[tlb.scala 41:26]
  reg [9:0] info_15; // @[tlb.scala 41:26]
  reg [31:0] pte_addr_0; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_1; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_2; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_3; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_4; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_5; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_6; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_7; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_8; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_9; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_10; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_11; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_12; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_13; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_14; // @[tlb.scala 42:30]
  reg [31:0] pte_addr_15; // @[tlb.scala 42:30]
  reg [1:0] pte_level_0; // @[tlb.scala 43:30]
  reg [1:0] pte_level_1; // @[tlb.scala 43:30]
  reg [1:0] pte_level_2; // @[tlb.scala 43:30]
  reg [1:0] pte_level_3; // @[tlb.scala 43:30]
  reg [1:0] pte_level_4; // @[tlb.scala 43:30]
  reg [1:0] pte_level_5; // @[tlb.scala 43:30]
  reg [1:0] pte_level_6; // @[tlb.scala 43:30]
  reg [1:0] pte_level_7; // @[tlb.scala 43:30]
  reg [1:0] pte_level_8; // @[tlb.scala 43:30]
  reg [1:0] pte_level_9; // @[tlb.scala 43:30]
  reg [1:0] pte_level_10; // @[tlb.scala 43:30]
  reg [1:0] pte_level_11; // @[tlb.scala 43:30]
  reg [1:0] pte_level_12; // @[tlb.scala 43:30]
  reg [1:0] pte_level_13; // @[tlb.scala 43:30]
  reg [1:0] pte_level_14; // @[tlb.scala 43:30]
  reg [1:0] pte_level_15; // @[tlb.scala 43:30]
  reg  valid_0; // @[tlb.scala 44:26]
  reg  valid_1; // @[tlb.scala 44:26]
  reg  valid_2; // @[tlb.scala 44:26]
  reg  valid_3; // @[tlb.scala 44:26]
  reg  valid_4; // @[tlb.scala 44:26]
  reg  valid_5; // @[tlb.scala 44:26]
  reg  valid_6; // @[tlb.scala 44:26]
  reg  valid_7; // @[tlb.scala 44:26]
  reg  valid_8; // @[tlb.scala 44:26]
  reg  valid_9; // @[tlb.scala 44:26]
  reg  valid_10; // @[tlb.scala 44:26]
  reg  valid_11; // @[tlb.scala 44:26]
  reg  valid_12; // @[tlb.scala 44:26]
  reg  valid_13; // @[tlb.scala 44:26]
  reg  valid_14; // @[tlb.scala 44:26]
  reg  valid_15; // @[tlb.scala 44:26]
  reg [63:0] pre_addr; // @[tlb.scala 46:30]
  reg [31:0] pte_addr_r; // @[tlb.scala 47:30]
  reg [63:0] wpte_data_r; // @[tlb.scala 48:30]
  reg [4:0] dc_mode_r; // @[tlb.scala 49:30]
  reg  out_valid_r; // @[tlb.scala 51:30]
  reg [31:0] out_paddr_r; // @[tlb.scala 52:30]
  reg [63:0] out_excep_r_cause; // @[tlb.scala 53:30]
  reg [63:0] out_excep_r_tval; // @[tlb.scala 53:30]
  reg  out_excep_r_en; // @[tlb.scala 53:30]
  wire [51:0] inp_tag = io_va2pa_vaddr[63:12]; // @[tlb.scala 58:33]
  wire  _mode_T = io_va2pa_m_type == 2'h1; // @[tlb.scala 61:26]
  wire [1:0] _mode_T_3 = io_mmuState_mstatus[17] ? io_mmuState_mstatus[12:11] : io_mmuState_priv; // @[Mux.scala 47:69]
  wire [1:0] mode = _mode_T ? io_mmuState_priv : _mode_T_3; // @[Mux.scala 47:69]
  wire [3:0] mmuMode = mode == 2'h3 ? 4'h0 : io_mmuState_satp[63:60]; // @[tlb.scala 65:22]
  wire  is_Sv39 = mmuMode == 4'h8; // @[tlb.scala 66:27]
  wire [51:0] _tlb_tag_mask_T_4 = 2'h0 == pte_level_0 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_6 = 2'h1 == pte_level_0 ? 52'hffffffffffe00 : _tlb_tag_mask_T_4; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask = 2'h2 == pte_level_0 ? 52'hffffffffc0000 : _tlb_tag_mask_T_6; // @[Mux.scala 80:57]
  wire [51:0] _T_1 = inp_tag & tlb_tag_mask; // @[tlb.scala 73:24]
  wire [19:0] _GEN_2 = _T_1 == tag_0 & valid_0 ? paddr_0 : 20'h0; // @[tlb.scala 73:64 tlb.scala 75:28 tlb.scala 68:40]
  wire [9:0] _GEN_4 = _T_1 == tag_0 & valid_0 ? info_0 : 10'h0; // @[tlb.scala 73:64 tlb.scala 77:28 tlb.scala 68:86]
  wire [31:0] _GEN_5 = _T_1 == tag_0 & valid_0 ? pte_addr_0 : 32'h0; // @[tlb.scala 73:64 tlb.scala 78:31 tlb.scala 69:23]
  wire [1:0] _GEN_7 = _T_1 == tag_0 & valid_0 ? pte_level_0 : 2'h0; // @[tlb.scala 73:64 tlb.scala 80:31 tlb.scala 69:69]
  wire [51:0] _tlb_tag_mask_T_12 = 2'h0 == pte_level_1 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_14 = 2'h1 == pte_level_1 ? 52'hffffffffffe00 : _tlb_tag_mask_T_12; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_1 = 2'h2 == pte_level_1 ? 52'hffffffffc0000 : _tlb_tag_mask_T_14; // @[Mux.scala 80:57]
  wire [51:0] _T_4 = inp_tag & tlb_tag_mask_1; // @[tlb.scala 73:24]
  wire  _T_6 = _T_4 == tag_1 & valid_1; // @[tlb.scala 73:52]
  wire [19:0] _GEN_9 = _T_4 == tag_1 & valid_1 ? paddr_1 : _GEN_2; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_11 = _T_4 == tag_1 & valid_1 ? info_1 : _GEN_4; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_12 = _T_4 == tag_1 & valid_1 ? pte_addr_1 : _GEN_5; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [1:0] _GEN_14 = _T_4 == tag_1 & valid_1 ? pte_level_1 : _GEN_7; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_20 = 2'h0 == pte_level_2 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_22 = 2'h1 == pte_level_2 ? 52'hffffffffffe00 : _tlb_tag_mask_T_20; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_2 = 2'h2 == pte_level_2 ? 52'hffffffffc0000 : _tlb_tag_mask_T_22; // @[Mux.scala 80:57]
  wire [51:0] _T_7 = inp_tag & tlb_tag_mask_2; // @[tlb.scala 73:24]
  wire [19:0] _GEN_16 = _T_7 == tag_2 & valid_2 ? paddr_2 : _GEN_9; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_18 = _T_7 == tag_2 & valid_2 ? info_2 : _GEN_11; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_19 = _T_7 == tag_2 & valid_2 ? pte_addr_2 : _GEN_12; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [1:0] _GEN_20 = _T_7 == tag_2 & valid_2 ? 2'h2 : {{1'd0}, _T_6}; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_21 = _T_7 == tag_2 & valid_2 ? pte_level_2 : _GEN_14; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_28 = 2'h0 == pte_level_3 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_30 = 2'h1 == pte_level_3 ? 52'hffffffffffe00 : _tlb_tag_mask_T_28; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_3 = 2'h2 == pte_level_3 ? 52'hffffffffc0000 : _tlb_tag_mask_T_30; // @[Mux.scala 80:57]
  wire [51:0] _T_10 = inp_tag & tlb_tag_mask_3; // @[tlb.scala 73:24]
  wire [19:0] _GEN_23 = _T_10 == tag_3 & valid_3 ? paddr_3 : _GEN_16; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_25 = _T_10 == tag_3 & valid_3 ? info_3 : _GEN_18; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_26 = _T_10 == tag_3 & valid_3 ? pte_addr_3 : _GEN_19; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [1:0] _GEN_27 = _T_10 == tag_3 & valid_3 ? 2'h3 : _GEN_20; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_28 = _T_10 == tag_3 & valid_3 ? pte_level_3 : _GEN_21; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_36 = 2'h0 == pte_level_4 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_38 = 2'h1 == pte_level_4 ? 52'hffffffffffe00 : _tlb_tag_mask_T_36; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_4 = 2'h2 == pte_level_4 ? 52'hffffffffc0000 : _tlb_tag_mask_T_38; // @[Mux.scala 80:57]
  wire [51:0] _T_13 = inp_tag & tlb_tag_mask_4; // @[tlb.scala 73:24]
  wire [19:0] _GEN_30 = _T_13 == tag_4 & valid_4 ? paddr_4 : _GEN_23; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_32 = _T_13 == tag_4 & valid_4 ? info_4 : _GEN_25; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_33 = _T_13 == tag_4 & valid_4 ? pte_addr_4 : _GEN_26; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [2:0] _GEN_34 = _T_13 == tag_4 & valid_4 ? 3'h4 : {{1'd0}, _GEN_27}; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_35 = _T_13 == tag_4 & valid_4 ? pte_level_4 : _GEN_28; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_44 = 2'h0 == pte_level_5 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_46 = 2'h1 == pte_level_5 ? 52'hffffffffffe00 : _tlb_tag_mask_T_44; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_5 = 2'h2 == pte_level_5 ? 52'hffffffffc0000 : _tlb_tag_mask_T_46; // @[Mux.scala 80:57]
  wire [51:0] _T_16 = inp_tag & tlb_tag_mask_5; // @[tlb.scala 73:24]
  wire [19:0] _GEN_37 = _T_16 == tag_5 & valid_5 ? paddr_5 : _GEN_30; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_39 = _T_16 == tag_5 & valid_5 ? info_5 : _GEN_32; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_40 = _T_16 == tag_5 & valid_5 ? pte_addr_5 : _GEN_33; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [2:0] _GEN_41 = _T_16 == tag_5 & valid_5 ? 3'h5 : _GEN_34; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_42 = _T_16 == tag_5 & valid_5 ? pte_level_5 : _GEN_35; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_52 = 2'h0 == pte_level_6 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_54 = 2'h1 == pte_level_6 ? 52'hffffffffffe00 : _tlb_tag_mask_T_52; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_6 = 2'h2 == pte_level_6 ? 52'hffffffffc0000 : _tlb_tag_mask_T_54; // @[Mux.scala 80:57]
  wire [51:0] _T_19 = inp_tag & tlb_tag_mask_6; // @[tlb.scala 73:24]
  wire [19:0] _GEN_44 = _T_19 == tag_6 & valid_6 ? paddr_6 : _GEN_37; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_46 = _T_19 == tag_6 & valid_6 ? info_6 : _GEN_39; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_47 = _T_19 == tag_6 & valid_6 ? pte_addr_6 : _GEN_40; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [2:0] _GEN_48 = _T_19 == tag_6 & valid_6 ? 3'h6 : _GEN_41; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_49 = _T_19 == tag_6 & valid_6 ? pte_level_6 : _GEN_42; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_60 = 2'h0 == pte_level_7 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_62 = 2'h1 == pte_level_7 ? 52'hffffffffffe00 : _tlb_tag_mask_T_60; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_7 = 2'h2 == pte_level_7 ? 52'hffffffffc0000 : _tlb_tag_mask_T_62; // @[Mux.scala 80:57]
  wire [51:0] _T_22 = inp_tag & tlb_tag_mask_7; // @[tlb.scala 73:24]
  wire [19:0] _GEN_51 = _T_22 == tag_7 & valid_7 ? paddr_7 : _GEN_44; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_53 = _T_22 == tag_7 & valid_7 ? info_7 : _GEN_46; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_54 = _T_22 == tag_7 & valid_7 ? pte_addr_7 : _GEN_47; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [2:0] _GEN_55 = _T_22 == tag_7 & valid_7 ? 3'h7 : _GEN_48; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_56 = _T_22 == tag_7 & valid_7 ? pte_level_7 : _GEN_49; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_68 = 2'h0 == pte_level_8 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_70 = 2'h1 == pte_level_8 ? 52'hffffffffffe00 : _tlb_tag_mask_T_68; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_8 = 2'h2 == pte_level_8 ? 52'hffffffffc0000 : _tlb_tag_mask_T_70; // @[Mux.scala 80:57]
  wire [51:0] _T_25 = inp_tag & tlb_tag_mask_8; // @[tlb.scala 73:24]
  wire [19:0] _GEN_58 = _T_25 == tag_8 & valid_8 ? paddr_8 : _GEN_51; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_60 = _T_25 == tag_8 & valid_8 ? info_8 : _GEN_53; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_61 = _T_25 == tag_8 & valid_8 ? pte_addr_8 : _GEN_54; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [3:0] _GEN_62 = _T_25 == tag_8 & valid_8 ? 4'h8 : {{1'd0}, _GEN_55}; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_63 = _T_25 == tag_8 & valid_8 ? pte_level_8 : _GEN_56; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_76 = 2'h0 == pte_level_9 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_78 = 2'h1 == pte_level_9 ? 52'hffffffffffe00 : _tlb_tag_mask_T_76; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_9 = 2'h2 == pte_level_9 ? 52'hffffffffc0000 : _tlb_tag_mask_T_78; // @[Mux.scala 80:57]
  wire [51:0] _T_28 = inp_tag & tlb_tag_mask_9; // @[tlb.scala 73:24]
  wire  _GEN_64 = _T_28 == tag_9 & valid_9 | (_T_25 == tag_8 & valid_8 | (_T_22 == tag_7 & valid_7 | (_T_19 == tag_6 &
    valid_6 | (_T_16 == tag_5 & valid_5 | (_T_13 == tag_4 & valid_4 | (_T_10 == tag_3 & valid_3 | (_T_7 == tag_2 &
    valid_2 | (_T_4 == tag_1 & valid_1 | _T_1 == tag_0 & valid_0)))))))); // @[tlb.scala 73:64 tlb.scala 74:28]
  wire [19:0] _GEN_65 = _T_28 == tag_9 & valid_9 ? paddr_9 : _GEN_58; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_67 = _T_28 == tag_9 & valid_9 ? info_9 : _GEN_60; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_68 = _T_28 == tag_9 & valid_9 ? pte_addr_9 : _GEN_61; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [3:0] _GEN_69 = _T_28 == tag_9 & valid_9 ? 4'h9 : _GEN_62; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_70 = _T_28 == tag_9 & valid_9 ? pte_level_9 : _GEN_63; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_84 = 2'h0 == pte_level_10 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_86 = 2'h1 == pte_level_10 ? 52'hffffffffffe00 : _tlb_tag_mask_T_84; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_10 = 2'h2 == pte_level_10 ? 52'hffffffffc0000 : _tlb_tag_mask_T_86; // @[Mux.scala 80:57]
  wire [51:0] _T_31 = inp_tag & tlb_tag_mask_10; // @[tlb.scala 73:24]
  wire [19:0] _GEN_72 = _T_31 == tag_10 & valid_10 ? paddr_10 : _GEN_65; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_74 = _T_31 == tag_10 & valid_10 ? info_10 : _GEN_67; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_75 = _T_31 == tag_10 & valid_10 ? pte_addr_10 : _GEN_68; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [3:0] _GEN_76 = _T_31 == tag_10 & valid_10 ? 4'ha : _GEN_69; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_77 = _T_31 == tag_10 & valid_10 ? pte_level_10 : _GEN_70; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_92 = 2'h0 == pte_level_11 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_94 = 2'h1 == pte_level_11 ? 52'hffffffffffe00 : _tlb_tag_mask_T_92; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_11 = 2'h2 == pte_level_11 ? 52'hffffffffc0000 : _tlb_tag_mask_T_94; // @[Mux.scala 80:57]
  wire [51:0] _T_34 = inp_tag & tlb_tag_mask_11; // @[tlb.scala 73:24]
  wire [19:0] _GEN_79 = _T_34 == tag_11 & valid_11 ? paddr_11 : _GEN_72; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_81 = _T_34 == tag_11 & valid_11 ? info_11 : _GEN_74; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_82 = _T_34 == tag_11 & valid_11 ? pte_addr_11 : _GEN_75; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [3:0] _GEN_83 = _T_34 == tag_11 & valid_11 ? 4'hb : _GEN_76; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_84 = _T_34 == tag_11 & valid_11 ? pte_level_11 : _GEN_77; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_100 = 2'h0 == pte_level_12 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_102 = 2'h1 == pte_level_12 ? 52'hffffffffffe00 : _tlb_tag_mask_T_100; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_12 = 2'h2 == pte_level_12 ? 52'hffffffffc0000 : _tlb_tag_mask_T_102; // @[Mux.scala 80:57]
  wire [51:0] _T_37 = inp_tag & tlb_tag_mask_12; // @[tlb.scala 73:24]
  wire [19:0] _GEN_86 = _T_37 == tag_12 & valid_12 ? paddr_12 : _GEN_79; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_88 = _T_37 == tag_12 & valid_12 ? info_12 : _GEN_81; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_89 = _T_37 == tag_12 & valid_12 ? pte_addr_12 : _GEN_82; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [3:0] _GEN_90 = _T_37 == tag_12 & valid_12 ? 4'hc : _GEN_83; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_91 = _T_37 == tag_12 & valid_12 ? pte_level_12 : _GEN_84; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_108 = 2'h0 == pte_level_13 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_110 = 2'h1 == pte_level_13 ? 52'hffffffffffe00 : _tlb_tag_mask_T_108; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_13 = 2'h2 == pte_level_13 ? 52'hffffffffc0000 : _tlb_tag_mask_T_110; // @[Mux.scala 80:57]
  wire [51:0] _T_40 = inp_tag & tlb_tag_mask_13; // @[tlb.scala 73:24]
  wire [19:0] _GEN_93 = _T_40 == tag_13 & valid_13 ? paddr_13 : _GEN_86; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_95 = _T_40 == tag_13 & valid_13 ? info_13 : _GEN_88; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_96 = _T_40 == tag_13 & valid_13 ? pte_addr_13 : _GEN_89; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [3:0] _GEN_97 = _T_40 == tag_13 & valid_13 ? 4'hd : _GEN_90; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_98 = _T_40 == tag_13 & valid_13 ? pte_level_13 : _GEN_91; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_116 = 2'h0 == pte_level_14 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_118 = 2'h1 == pte_level_14 ? 52'hffffffffffe00 : _tlb_tag_mask_T_116; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_14 = 2'h2 == pte_level_14 ? 52'hffffffffc0000 : _tlb_tag_mask_T_118; // @[Mux.scala 80:57]
  wire [51:0] _T_43 = inp_tag & tlb_tag_mask_14; // @[tlb.scala 73:24]
  wire [19:0] _GEN_100 = _T_43 == tag_14 & valid_14 ? paddr_14 : _GEN_93; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] _GEN_102 = _T_43 == tag_14 & valid_14 ? info_14 : _GEN_95; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] _GEN_103 = _T_43 == tag_14 & valid_14 ? pte_addr_14 : _GEN_96; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [3:0] _GEN_104 = _T_43 == tag_14 & valid_14 ? 4'he : _GEN_97; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] _GEN_105 = _T_43 == tag_14 & valid_14 ? pte_level_14 : _GEN_98; // @[tlb.scala 73:64 tlb.scala 80:31]
  wire [51:0] _tlb_tag_mask_T_124 = 2'h0 == pte_level_15 ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _tlb_tag_mask_T_126 = 2'h1 == pte_level_15 ? 52'hffffffffffe00 : _tlb_tag_mask_T_124; // @[Mux.scala 80:57]
  wire [51:0] tlb_tag_mask_15 = 2'h2 == pte_level_15 ? 52'hffffffffc0000 : _tlb_tag_mask_T_126; // @[Mux.scala 80:57]
  wire [51:0] _T_46 = inp_tag & tlb_tag_mask_15; // @[tlb.scala 73:24]
  wire  tlbMsg_tlbHit = _T_46 == tag_15 & valid_15 | (_T_43 == tag_14 & valid_14 | (_T_40 == tag_13 & valid_13 | (_T_37
     == tag_12 & valid_12 | (_T_34 == tag_11 & valid_11 | (_T_31 == tag_10 & valid_10 | _GEN_64))))); // @[tlb.scala 73:64 tlb.scala 74:28]
  wire [19:0] tlbMsg_tlbPa = _T_46 == tag_15 & valid_15 ? paddr_15 : _GEN_100; // @[tlb.scala 73:64 tlb.scala 75:28]
  wire [9:0] tlbMsg_tlbInfo = _T_46 == tag_15 & valid_15 ? info_15 : _GEN_102; // @[tlb.scala 73:64 tlb.scala 77:28]
  wire [31:0] tlbMsg_tlbPteAddr = _T_46 == tag_15 & valid_15 ? pte_addr_15 : _GEN_103; // @[tlb.scala 73:64 tlb.scala 78:31]
  wire [3:0] tlbMsg_tlbIdx = _T_46 == tag_15 & valid_15 ? 4'hf : _GEN_104; // @[tlb.scala 73:64 tlb.scala 79:28]
  wire [1:0] tlbMsg_tlbLevel = _T_46 == tag_15 & valid_15 ? pte_level_15 : _GEN_105; // @[tlb.scala 73:64 tlb.scala 80:31]
  reg [1:0] state; // @[tlb.scala 84:24]
  reg  flush_r; // @[tlb.scala 85:26]
  wire  _T_50 = state == 2'h0; // @[tlb.scala 87:20]
  wire  _GEN_113 = state == 2'h0 ? 1'h0 : valid_0; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_114 = state == 2'h0 ? 1'h0 : valid_1; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_115 = state == 2'h0 ? 1'h0 : valid_2; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_116 = state == 2'h0 ? 1'h0 : valid_3; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_117 = state == 2'h0 ? 1'h0 : valid_4; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_118 = state == 2'h0 ? 1'h0 : valid_5; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_119 = state == 2'h0 ? 1'h0 : valid_6; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_120 = state == 2'h0 ? 1'h0 : valid_7; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_121 = state == 2'h0 ? 1'h0 : valid_8; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_122 = state == 2'h0 ? 1'h0 : valid_9; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_123 = state == 2'h0 ? 1'h0 : valid_10; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_124 = state == 2'h0 ? 1'h0 : valid_11; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_125 = state == 2'h0 ? 1'h0 : valid_12; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_126 = state == 2'h0 ? 1'h0 : valid_13; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_127 = state == 2'h0 ? 1'h0 : valid_14; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_128 = state == 2'h0 ? 1'h0 : valid_15; // @[tlb.scala 87:30 tlb.scala 88:19 tlb.scala 44:26]
  wire  _GEN_130 = io_flush | flush_r ? _GEN_113 : valid_0; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_131 = io_flush | flush_r ? _GEN_114 : valid_1; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_132 = io_flush | flush_r ? _GEN_115 : valid_2; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_133 = io_flush | flush_r ? _GEN_116 : valid_3; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_134 = io_flush | flush_r ? _GEN_117 : valid_4; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_135 = io_flush | flush_r ? _GEN_118 : valid_5; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_136 = io_flush | flush_r ? _GEN_119 : valid_6; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_137 = io_flush | flush_r ? _GEN_120 : valid_7; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_138 = io_flush | flush_r ? _GEN_121 : valid_8; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_139 = io_flush | flush_r ? _GEN_122 : valid_9; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_140 = io_flush | flush_r ? _GEN_123 : valid_10; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_141 = io_flush | flush_r ? _GEN_124 : valid_11; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_142 = io_flush | flush_r ? _GEN_125 : valid_12; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_143 = io_flush | flush_r ? _GEN_126 : valid_13; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_144 = io_flush | flush_r ? _GEN_127 : valid_14; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  _GEN_145 = io_flush | flush_r ? _GEN_128 : valid_15; // @[tlb.scala 86:30 tlb.scala 44:26]
  wire  handshake = io_va2pa_vvalid & io_va2pa_ready; // @[tlb.scala 94:37]
  reg [1:0] m_type_r; // @[tlb.scala 95:27]
  wire [1:0] cur_m_type = handshake ? io_va2pa_m_type : m_type_r; // @[tlb.scala 96:25]
  wire  _ad_T = cur_m_type == 2'h3; // @[common.scala 243:20]
  wire [9:0] ad = cur_m_type == 2'h3 ? 10'hc0 : 10'h40; // @[common.scala 243:12]
  wire  _GEN_150 = io_va2pa_pvalid | io_va2pa_tlb_excep_en ? 1'h0 : out_valid_r; // @[tlb.scala 108:51 tlb.scala 109:21 tlb.scala 51:30]
  wire  _GEN_151 = io_va2pa_pvalid | io_va2pa_tlb_excep_en ? 1'h0 : out_excep_r_en; // @[tlb.scala 108:51 tlb.scala 110:24 tlb.scala 53:30]
  wire  dc_hand = io_dcacheRW_ready & io_dcacheRW_dc_mode != 5'h0; // @[tlb.scala 122:37]
  wire [24:0] _tlb_high_legal_T_2 = io_va2pa_vaddr[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire  tlb_high_legal = _tlb_high_legal_T_2 == io_va2pa_vaddr[63:39]; // @[tlb.scala 125:55]
  wire  _tlb_access_illegal_T_11 = cur_m_type == 2'h2 & ~(tlbMsg_tlbInfo[1] | io_mmuState_mstatus[19] & tlbMsg_tlbInfo[3
    ]); // @[tlb.scala 127:60]
  wire  _tlb_access_illegal_T_12 = cur_m_type == 2'h1 & ~tlbMsg_tlbInfo[3] | _tlb_access_illegal_T_11; // @[tlb.scala 126:89]
  wire  _tlb_access_illegal_T_16 = _ad_T & ~tlbMsg_tlbInfo[2]; // @[tlb.scala 128:57]
  wire  tlb_access_illegal = _tlb_access_illegal_T_12 | _tlb_access_illegal_T_16; // @[tlb.scala 127:152]
  wire [3:0] select = {select_prng_io_out_3,select_prng_io_out_2,select_prng_io_out_1,select_prng_io_out_0}; // @[PRNG.scala 86:17]
  reg [3:0] select_r; // @[tlb.scala 130:27]
  reg [7:0] offset; // @[tlb.scala 131:26]
  reg [1:0] level; // @[tlb.scala 132:26]
  reg  wpte_hs_r; // @[tlb.scala 134:28]
  wire  _T_54 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire [63:0] _out_excep_r_cause_T_1 = 2'h1 == io_va2pa_m_type ? 64'hc : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _out_excep_r_cause_T_3 = 2'h2 == io_va2pa_m_type ? 64'hd : _out_excep_r_cause_T_1; // @[Mux.scala 80:57]
  wire [63:0] _out_excep_r_cause_T_5 = 2'h3 == io_va2pa_m_type ? 64'hf : _out_excep_r_cause_T_3; // @[Mux.scala 80:57]
  wire [51:0] _paddr_mask_T_4 = 2'h0 == tlbMsg_tlbLevel ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _paddr_mask_T_6 = 2'h1 == tlbMsg_tlbLevel ? 52'hffffffffffe00 : _paddr_mask_T_4; // @[Mux.scala 80:57]
  wire [51:0] paddr_mask_hi = 2'h2 == tlbMsg_tlbLevel ? 52'hffffffffc0000 : _paddr_mask_T_6; // @[Mux.scala 80:57]
  wire [63:0] paddr_mask = {paddr_mask_hi,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _out_paddr_r_T = {tlbMsg_tlbPa, 12'h0}; // @[tlb.scala 148:93]
  wire [63:0] _out_paddr_r_T_1 = ~paddr_mask; // @[common.scala 201:19]
  wire [63:0] _out_paddr_r_T_2 = io_va2pa_vaddr & _out_paddr_r_T_1; // @[common.scala 201:17]
  wire [63:0] _GEN_1417 = {{32'd0}, _out_paddr_r_T}; // @[common.scala 201:36]
  wire [63:0] _out_paddr_r_T_3 = _GEN_1417 & paddr_mask; // @[common.scala 201:36]
  wire [63:0] _out_paddr_r_T_4 = _out_paddr_r_T_2 | _out_paddr_r_T_3; // @[common.scala 201:26]
  wire [9:0] _T_59 = ad & tlbMsg_tlbInfo; // @[tlb.scala 149:30]
  wire [9:0] wpte_data_r_lo = tlbMsg_tlbInfo | ad; // @[tlb.scala 153:84]
  wire [63:0] _wpte_data_r_T = {34'h0,tlbMsg_tlbPa,wpte_data_r_lo}; // @[Cat.scala 30:58]
  wire [9:0] _GEN_152 = 4'h0 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_0; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_153 = 4'h1 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_1; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_154 = 4'h2 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_2; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_155 = 4'h3 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_3; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_156 = 4'h4 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_4; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_157 = 4'h5 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_5; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_158 = 4'h6 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_6; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_159 = 4'h7 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_7; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_160 = 4'h8 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_8; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_161 = 4'h9 == tlbMsg_tlbIdx ? wpte_data_r_lo : info_9; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_162 = 4'ha == tlbMsg_tlbIdx ? wpte_data_r_lo : info_10; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_163 = 4'hb == tlbMsg_tlbIdx ? wpte_data_r_lo : info_11; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_164 = 4'hc == tlbMsg_tlbIdx ? wpte_data_r_lo : info_12; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_165 = 4'hd == tlbMsg_tlbIdx ? wpte_data_r_lo : info_13; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_166 = 4'he == tlbMsg_tlbIdx ? wpte_data_r_lo : info_14; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [9:0] _GEN_167 = 4'hf == tlbMsg_tlbIdx ? wpte_data_r_lo : info_15; // @[tlb.scala 154:45 tlb.scala 154:45 tlb.scala 41:26]
  wire [1:0] _GEN_168 = _T_59 != ad & is_Sv39 ? 2'h3 : state; // @[tlb.scala 149:66 tlb.scala 150:31 tlb.scala 84:24]
  wire  _GEN_169 = _T_59 != ad & is_Sv39 ? 1'h0 : wpte_hs_r; // @[tlb.scala 149:66 tlb.scala 151:35 tlb.scala 134:28]
  wire [31:0] _GEN_170 = _T_59 != ad & is_Sv39 ? tlbMsg_tlbPteAddr : pte_addr_r; // @[tlb.scala 149:66 tlb.scala 152:37 tlb.scala 47:30]
  wire [63:0] _GEN_171 = _T_59 != ad & is_Sv39 ? _wpte_data_r_T : wpte_data_r; // @[tlb.scala 149:66 tlb.scala 153:37 tlb.scala 48:30]
  wire [9:0] _GEN_172 = _T_59 != ad & is_Sv39 ? _GEN_152 : info_0; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_173 = _T_59 != ad & is_Sv39 ? _GEN_153 : info_1; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_174 = _T_59 != ad & is_Sv39 ? _GEN_154 : info_2; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_175 = _T_59 != ad & is_Sv39 ? _GEN_155 : info_3; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_176 = _T_59 != ad & is_Sv39 ? _GEN_156 : info_4; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_177 = _T_59 != ad & is_Sv39 ? _GEN_157 : info_5; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_178 = _T_59 != ad & is_Sv39 ? _GEN_158 : info_6; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_179 = _T_59 != ad & is_Sv39 ? _GEN_159 : info_7; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_180 = _T_59 != ad & is_Sv39 ? _GEN_160 : info_8; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_181 = _T_59 != ad & is_Sv39 ? _GEN_161 : info_9; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_182 = _T_59 != ad & is_Sv39 ? _GEN_162 : info_10; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_183 = _T_59 != ad & is_Sv39 ? _GEN_163 : info_11; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_184 = _T_59 != ad & is_Sv39 ? _GEN_164 : info_12; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_185 = _T_59 != ad & is_Sv39 ? _GEN_165 : info_13; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_186 = _T_59 != ad & is_Sv39 ? _GEN_166 : info_14; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [9:0] _GEN_187 = _T_59 != ad & is_Sv39 ? _GEN_167 : info_15; // @[tlb.scala 149:66 tlb.scala 41:26]
  wire [43:0] pte_addr_r_hi_hi = io_mmuState_satp[43:0]; // @[tlb.scala 166:59]
  wire [63:0] _pte_addr_r_T = {{30'd0}, io_va2pa_vaddr[63:30]}; // @[tlb.scala 166:83]
  wire [8:0] pte_addr_r_hi_lo = _pte_addr_r_T[8:0]; // @[tlb.scala 166:91]
  wire [55:0] _pte_addr_r_T_1 = {pte_addr_r_hi_hi,pte_addr_r_hi_lo,3'h0}; // @[Cat.scala 30:58]
  wire  _GEN_188 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 | _GEN_151; // @[tlb.scala 162:81 tlb.scala 164:40]
  wire [55:0] _GEN_189 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 ? {{24'd0}, pte_addr_r} : _pte_addr_r_T_1; // @[tlb.scala 162:81 tlb.scala 47:30 tlb.scala 166:36]
  wire [4:0] _GEN_190 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 ? 5'h0 : 5'h7; // @[tlb.scala 162:81 tlb.scala 138:27 tlb.scala 167:36]
  wire [7:0] _GEN_191 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 ? offset : 8'h1e; // @[tlb.scala 162:81 tlb.scala 131:26 tlb.scala 168:33]
  wire [1:0] _GEN_192 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 ? level : 2'h3; // @[tlb.scala 162:81 tlb.scala 132:26 tlb.scala 169:33]
  wire [1:0] _GEN_194 = ~tlbMsg_tlbHit ? 2'h1 : state; // @[tlb.scala 156:43 tlb.scala 84:24]
  wire [3:0] _GEN_195 = ~tlbMsg_tlbHit ? select : select_r; // @[tlb.scala 156:43 tlb.scala 158:32 tlb.scala 130:27]
  wire [1:0] _GEN_196 = ~tlbMsg_tlbHit ? io_va2pa_m_type : m_type_r; // @[tlb.scala 156:43 tlb.scala 159:32 tlb.scala 95:27]
  wire [63:0] _GEN_197 = ~tlbMsg_tlbHit ? _out_excep_r_cause_T_5 : out_excep_r_cause; // @[tlb.scala 156:43 tlb.scala 160:39 tlb.scala 53:30]
  wire [63:0] _GEN_198 = ~tlbMsg_tlbHit ? io_va2pa_vaddr : out_excep_r_tval; // @[tlb.scala 156:43 tlb.scala 161:39 tlb.scala 53:30]
  wire  _GEN_199 = ~tlbMsg_tlbHit ? _GEN_188 : _GEN_151; // @[tlb.scala 156:43]
  wire [55:0] _GEN_200 = ~tlbMsg_tlbHit ? _GEN_189 : {{24'd0}, pte_addr_r}; // @[tlb.scala 156:43 tlb.scala 47:30]
  wire [4:0] _GEN_201 = ~tlbMsg_tlbHit ? _GEN_190 : 5'h0; // @[tlb.scala 156:43 tlb.scala 138:27]
  wire [7:0] _GEN_202 = ~tlbMsg_tlbHit ? _GEN_191 : offset; // @[tlb.scala 156:43 tlb.scala 131:26]
  wire [1:0] _GEN_203 = ~tlbMsg_tlbHit ? _GEN_192 : level; // @[tlb.scala 156:43 tlb.scala 132:26]
  wire  _GEN_204 = tlbMsg_tlbHit | _GEN_150; // @[tlb.scala 144:42 tlb.scala 145:33]
  wire [63:0] _GEN_205 = tlbMsg_tlbHit ? _out_paddr_r_T_4 : {{32'd0}, out_paddr_r}; // @[tlb.scala 144:42 tlb.scala 148:33 tlb.scala 52:30]
  wire [1:0] _GEN_206 = tlbMsg_tlbHit ? _GEN_168 : _GEN_194; // @[tlb.scala 144:42]
  wire  _GEN_207 = tlbMsg_tlbHit ? _GEN_169 : wpte_hs_r; // @[tlb.scala 144:42 tlb.scala 134:28]
  wire [55:0] _GEN_208 = tlbMsg_tlbHit ? {{24'd0}, _GEN_170} : _GEN_200; // @[tlb.scala 144:42]
  wire [63:0] _GEN_209 = tlbMsg_tlbHit ? _GEN_171 : wpte_data_r; // @[tlb.scala 144:42 tlb.scala 48:30]
  wire [9:0] _GEN_210 = tlbMsg_tlbHit ? _GEN_172 : info_0; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_211 = tlbMsg_tlbHit ? _GEN_173 : info_1; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_212 = tlbMsg_tlbHit ? _GEN_174 : info_2; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_213 = tlbMsg_tlbHit ? _GEN_175 : info_3; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_214 = tlbMsg_tlbHit ? _GEN_176 : info_4; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_215 = tlbMsg_tlbHit ? _GEN_177 : info_5; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_216 = tlbMsg_tlbHit ? _GEN_178 : info_6; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_217 = tlbMsg_tlbHit ? _GEN_179 : info_7; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_218 = tlbMsg_tlbHit ? _GEN_180 : info_8; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_219 = tlbMsg_tlbHit ? _GEN_181 : info_9; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_220 = tlbMsg_tlbHit ? _GEN_182 : info_10; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_221 = tlbMsg_tlbHit ? _GEN_183 : info_11; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_222 = tlbMsg_tlbHit ? _GEN_184 : info_12; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_223 = tlbMsg_tlbHit ? _GEN_185 : info_13; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_224 = tlbMsg_tlbHit ? _GEN_186 : info_14; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [9:0] _GEN_225 = tlbMsg_tlbHit ? _GEN_187 : info_15; // @[tlb.scala 144:42 tlb.scala 41:26]
  wire [3:0] _GEN_226 = tlbMsg_tlbHit ? select_r : _GEN_195; // @[tlb.scala 144:42 tlb.scala 130:27]
  wire [1:0] _GEN_227 = tlbMsg_tlbHit ? m_type_r : _GEN_196; // @[tlb.scala 144:42 tlb.scala 95:27]
  wire [63:0] _GEN_228 = tlbMsg_tlbHit ? out_excep_r_cause : _GEN_197; // @[tlb.scala 144:42 tlb.scala 53:30]
  wire [63:0] _GEN_229 = tlbMsg_tlbHit ? out_excep_r_tval : _GEN_198; // @[tlb.scala 144:42 tlb.scala 53:30]
  wire  _GEN_230 = tlbMsg_tlbHit ? _GEN_151 : _GEN_199; // @[tlb.scala 144:42]
  wire [4:0] _GEN_231 = tlbMsg_tlbHit ? 5'h0 : _GEN_201; // @[tlb.scala 144:42 tlb.scala 138:27]
  wire [7:0] _GEN_232 = tlbMsg_tlbHit ? offset : _GEN_202; // @[tlb.scala 144:42 tlb.scala 131:26]
  wire [1:0] _GEN_233 = tlbMsg_tlbHit ? level : _GEN_203; // @[tlb.scala 144:42 tlb.scala 132:26]
  wire  _GEN_234 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal | _GEN_230; // @[tlb.scala 140:85 tlb.scala 141:36]
  wire [63:0] _GEN_235 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? _out_excep_r_cause_T_5 : _GEN_228; // @[tlb.scala 140:85 tlb.scala 142:39]
  wire [63:0] _GEN_236 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? io_va2pa_vaddr : _GEN_229; // @[tlb.scala 140:85 tlb.scala 143:39]
  wire  _GEN_237 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? _GEN_150 : _GEN_204; // @[tlb.scala 140:85]
  wire [63:0] _GEN_238 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? {{32'd0}, out_paddr_r} : _GEN_205; // @[tlb.scala 140:85 tlb.scala 52:30]
  wire [1:0] _GEN_239 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? state : _GEN_206; // @[tlb.scala 140:85 tlb.scala 84:24]
  wire  _GEN_240 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? wpte_hs_r : _GEN_207; // @[tlb.scala 140:85 tlb.scala 134:28]
  wire [55:0] _GEN_241 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? {{24'd0}, pte_addr_r} : _GEN_208; // @[tlb.scala 140:85 tlb.scala 47:30]
  wire [63:0] _GEN_242 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? wpte_data_r : _GEN_209; // @[tlb.scala 140:85 tlb.scala 48:30]
  wire [9:0] _GEN_243 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_0 : _GEN_210; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_244 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_1 : _GEN_211; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_245 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_2 : _GEN_212; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_246 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_3 : _GEN_213; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_247 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_4 : _GEN_214; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_248 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_5 : _GEN_215; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_249 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_6 : _GEN_216; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_250 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_7 : _GEN_217; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_251 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_8 : _GEN_218; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_252 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_9 : _GEN_219; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_253 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_10 : _GEN_220; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_254 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_11 : _GEN_221; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_255 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_12 : _GEN_222; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_256 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_13 : _GEN_223; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_257 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_14 : _GEN_224; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [9:0] _GEN_258 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_15 : _GEN_225; // @[tlb.scala 140:85 tlb.scala 41:26]
  wire [3:0] _GEN_259 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? select_r : _GEN_226; // @[tlb.scala 140:85 tlb.scala 130:27]
  wire [1:0] _GEN_260 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? m_type_r : _GEN_227; // @[tlb.scala 140:85 tlb.scala 95:27]
  wire [4:0] _GEN_261 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? 5'h0 : _GEN_231; // @[tlb.scala 140:85 tlb.scala 138:27]
  wire [7:0] _GEN_262 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? offset : _GEN_232; // @[tlb.scala 140:85 tlb.scala 131:26]
  wire [1:0] _GEN_263 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? level : _GEN_233; // @[tlb.scala 140:85 tlb.scala 132:26]
  wire [63:0] _GEN_268 = ~handshake ? {{32'd0}, out_paddr_r} : _GEN_238; // @[tlb.scala 139:33 tlb.scala 52:30]
  wire [55:0] _GEN_271 = ~handshake ? {{24'd0}, pte_addr_r} : _GEN_241; // @[tlb.scala 139:33 tlb.scala 47:30]
  wire  _T_68 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [4:0] _dc_mode_r_T = wpte_hs_r ? 5'h0 : 5'hb; // @[tlb.scala 175:33]
  wire [4:0] _GEN_294 = io_dcacheRW_ready ? 5'h0 : _dc_mode_r_T; // @[tlb.scala 176:40 tlb.scala 177:31 tlb.scala 175:27]
  wire  _GEN_295 = io_dcacheRW_ready | wpte_hs_r; // @[tlb.scala 176:40 tlb.scala 178:31 tlb.scala 134:28]
  wire [1:0] _GEN_296 = io_dcacheRW_rvalid ? 2'h0 : state; // @[tlb.scala 180:41 tlb.scala 181:27 tlb.scala 84:24]
  wire  _T_69 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire [7:0] _offset_T_1 = offset - 8'h9; // @[tlb.scala 187:39]
  wire [1:0] _level_T_1 = level - 2'h1; // @[tlb.scala 188:38]
  wire [4:0] _GEN_297 = dc_hand ? 5'h0 : dc_mode_r; // @[tlb.scala 185:30 tlb.scala 186:31 tlb.scala 49:30]
  wire [7:0] _GEN_298 = dc_hand ? _offset_T_1 : offset; // @[tlb.scala 185:30 tlb.scala 187:29 tlb.scala 131:26]
  wire [1:0] _GEN_299 = dc_hand ? _level_T_1 : level; // @[tlb.scala 185:30 tlb.scala 188:29 tlb.scala 132:26]
  wire [63:0] _T_73 = io_dcacheRW_rdata & 64'hf; // @[tlb.scala 191:31]
  wire [63:0] _T_77 = io_dcacheRW_rdata & 64'hd0; // @[tlb.scala 192:35]
  wire [43:0] pte_addr_r_hi_hi_1 = io_dcacheRW_rdata[53:10]; // @[tlb.scala 196:50]
  wire [63:0] _pte_addr_r_T_2 = pre_addr >> offset; // @[tlb.scala 196:69]
  wire [8:0] pte_addr_r_hi_lo_1 = _pte_addr_r_T_2[8:0]; // @[tlb.scala 196:79]
  wire [55:0] _pte_addr_r_T_3 = {pte_addr_r_hi_hi_1,pte_addr_r_hi_lo_1,3'h0}; // @[Cat.scala 30:58]
  wire [1:0] _GEN_300 = _T_77 != 64'h0 ? 2'h0 : state; // @[tlb.scala 192:70 tlb.scala 193:35 tlb.scala 84:24]
  wire  _GEN_301 = _T_77 != 64'h0 | _GEN_151; // @[tlb.scala 192:70 tlb.scala 194:44]
  wire [55:0] _GEN_302 = _T_77 != 64'h0 ? {{24'd0}, pte_addr_r} : _pte_addr_r_T_3; // @[tlb.scala 192:70 tlb.scala 47:30 tlb.scala 196:40]
  wire [4:0] _GEN_303 = _T_77 != 64'h0 ? _GEN_297 : 5'h7; // @[tlb.scala 192:70 tlb.scala 197:40]
  wire  _T_83 = out_excep_r_cause == 64'hc; // @[tlb.scala 199:133]
  wire  _T_87 = io_dcacheRW_rdata[4] ? io_mmuState_priv == 2'h1 & (~io_mmuState_mstatus[18] | out_excep_r_cause == 64'hc
    ) : io_mmuState_priv == 2'h0; // @[tlb.scala 199:35]
  wire  _T_106 = out_excep_r_cause == 64'hd & ~(io_dcacheRW_rdata[1] | io_mmuState_mstatus[19] & io_dcacheRW_rdata[3]); // @[tlb.scala 208:82]
  wire  _T_107 = _T_83 & ~io_dcacheRW_rdata[3] | _T_106; // @[tlb.scala 207:102]
  wire  _T_111 = out_excep_r_cause == 64'hf & ~io_dcacheRW_rdata[2]; // @[tlb.scala 209:79]
  wire  _T_112 = _T_107 | _T_111; // @[tlb.scala 208:152]
  wire [51:0] _ppn_mask_T_4 = 2'h0 == level ? 52'hfffffffffffff : 52'h0; // @[Mux.scala 80:57]
  wire [51:0] _ppn_mask_T_6 = 2'h1 == level ? 52'hffffffffffe00 : _ppn_mask_T_4; // @[Mux.scala 80:57]
  wire [51:0] ppn_mask = 2'h2 == level ? 52'hffffffffc0000 : _ppn_mask_T_6; // @[Mux.scala 80:57]
  wire [51:0] _tag_T_1 = pre_addr[63:12] & ppn_mask; // @[tlb.scala 220:78]
  wire [51:0] _GEN_304 = 4'h0 == select_r ? _tag_T_1 : tag_0; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_305 = 4'h1 == select_r ? _tag_T_1 : tag_1; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_306 = 4'h2 == select_r ? _tag_T_1 : tag_2; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_307 = 4'h3 == select_r ? _tag_T_1 : tag_3; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_308 = 4'h4 == select_r ? _tag_T_1 : tag_4; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_309 = 4'h5 == select_r ? _tag_T_1 : tag_5; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_310 = 4'h6 == select_r ? _tag_T_1 : tag_6; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_311 = 4'h7 == select_r ? _tag_T_1 : tag_7; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_312 = 4'h8 == select_r ? _tag_T_1 : tag_8; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_313 = 4'h9 == select_r ? _tag_T_1 : tag_9; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_314 = 4'ha == select_r ? _tag_T_1 : tag_10; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_315 = 4'hb == select_r ? _tag_T_1 : tag_11; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_316 = 4'hc == select_r ? _tag_T_1 : tag_12; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_317 = 4'hd == select_r ? _tag_T_1 : tag_13; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_318 = 4'he == select_r ? _tag_T_1 : tag_14; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire [51:0] _GEN_319 = 4'hf == select_r ? _tag_T_1 : tag_15; // @[tlb.scala 220:39 tlb.scala 220:39 tlb.scala 39:26]
  wire  _GEN_320 = 4'h0 == select_r | _GEN_130; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_321 = 4'h1 == select_r | _GEN_131; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_322 = 4'h2 == select_r | _GEN_132; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_323 = 4'h3 == select_r | _GEN_133; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_324 = 4'h4 == select_r | _GEN_134; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_325 = 4'h5 == select_r | _GEN_135; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_326 = 4'h6 == select_r | _GEN_136; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_327 = 4'h7 == select_r | _GEN_137; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_328 = 4'h8 == select_r | _GEN_138; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_329 = 4'h9 == select_r | _GEN_139; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_330 = 4'ha == select_r | _GEN_140; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_331 = 4'hb == select_r | _GEN_141; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_332 = 4'hc == select_r | _GEN_142; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_333 = 4'hd == select_r | _GEN_143; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_334 = 4'he == select_r | _GEN_144; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire  _GEN_335 = 4'hf == select_r | _GEN_145; // @[tlb.scala 221:41 tlb.scala 221:41]
  wire [51:0] _GEN_1435 = {{32'd0}, io_dcacheRW_rdata[29:10]}; // @[tlb.scala 222:53]
  wire [51:0] update_pa = _GEN_1435 & ppn_mask; // @[tlb.scala 222:53]
  wire [19:0] _GEN_336 = 4'h0 == select_r ? update_pa[19:0] : paddr_0; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_337 = 4'h1 == select_r ? update_pa[19:0] : paddr_1; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_338 = 4'h2 == select_r ? update_pa[19:0] : paddr_2; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_339 = 4'h3 == select_r ? update_pa[19:0] : paddr_3; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_340 = 4'h4 == select_r ? update_pa[19:0] : paddr_4; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_341 = 4'h5 == select_r ? update_pa[19:0] : paddr_5; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_342 = 4'h6 == select_r ? update_pa[19:0] : paddr_6; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_343 = 4'h7 == select_r ? update_pa[19:0] : paddr_7; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_344 = 4'h8 == select_r ? update_pa[19:0] : paddr_8; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_345 = 4'h9 == select_r ? update_pa[19:0] : paddr_9; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_346 = 4'ha == select_r ? update_pa[19:0] : paddr_10; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_347 = 4'hb == select_r ? update_pa[19:0] : paddr_11; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_348 = 4'hc == select_r ? update_pa[19:0] : paddr_12; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_349 = 4'hd == select_r ? update_pa[19:0] : paddr_13; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_350 = 4'he == select_r ? update_pa[19:0] : paddr_14; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [19:0] _GEN_351 = 4'hf == select_r ? update_pa[19:0] : paddr_15; // @[tlb.scala 223:41 tlb.scala 223:41 tlb.scala 40:26]
  wire [31:0] _GEN_352 = 4'h0 == select_r ? pte_addr_r : pte_addr_0; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_353 = 4'h1 == select_r ? pte_addr_r : pte_addr_1; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_354 = 4'h2 == select_r ? pte_addr_r : pte_addr_2; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_355 = 4'h3 == select_r ? pte_addr_r : pte_addr_3; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_356 = 4'h4 == select_r ? pte_addr_r : pte_addr_4; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_357 = 4'h5 == select_r ? pte_addr_r : pte_addr_5; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_358 = 4'h6 == select_r ? pte_addr_r : pte_addr_6; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_359 = 4'h7 == select_r ? pte_addr_r : pte_addr_7; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_360 = 4'h8 == select_r ? pte_addr_r : pte_addr_8; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_361 = 4'h9 == select_r ? pte_addr_r : pte_addr_9; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_362 = 4'ha == select_r ? pte_addr_r : pte_addr_10; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_363 = 4'hb == select_r ? pte_addr_r : pte_addr_11; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_364 = 4'hc == select_r ? pte_addr_r : pte_addr_12; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_365 = 4'hd == select_r ? pte_addr_r : pte_addr_13; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_366 = 4'he == select_r ? pte_addr_r : pte_addr_14; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [31:0] _GEN_367 = 4'hf == select_r ? pte_addr_r : pte_addr_15; // @[tlb.scala 224:44 tlb.scala 224:44 tlb.scala 42:30]
  wire [1:0] _GEN_368 = 4'h0 == select_r ? level : pte_level_0; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_369 = 4'h1 == select_r ? level : pte_level_1; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_370 = 4'h2 == select_r ? level : pte_level_2; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_371 = 4'h3 == select_r ? level : pte_level_3; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_372 = 4'h4 == select_r ? level : pte_level_4; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_373 = 4'h5 == select_r ? level : pte_level_5; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_374 = 4'h6 == select_r ? level : pte_level_6; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_375 = 4'h7 == select_r ? level : pte_level_7; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_376 = 4'h8 == select_r ? level : pte_level_8; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_377 = 4'h9 == select_r ? level : pte_level_9; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_378 = 4'ha == select_r ? level : pte_level_10; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_379 = 4'hb == select_r ? level : pte_level_11; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_380 = 4'hc == select_r ? level : pte_level_12; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_381 = 4'hd == select_r ? level : pte_level_13; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_382 = 4'he == select_r ? level : pte_level_14; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [1:0] _GEN_383 = 4'hf == select_r ? level : pte_level_15; // @[tlb.scala 225:45 tlb.scala 225:45 tlb.scala 43:30]
  wire [9:0] _GEN_384 = 4'h0 == select_r ? io_dcacheRW_rdata[9:0] : info_0; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_385 = 4'h1 == select_r ? io_dcacheRW_rdata[9:0] : info_1; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_386 = 4'h2 == select_r ? io_dcacheRW_rdata[9:0] : info_2; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_387 = 4'h3 == select_r ? io_dcacheRW_rdata[9:0] : info_3; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_388 = 4'h4 == select_r ? io_dcacheRW_rdata[9:0] : info_4; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_389 = 4'h5 == select_r ? io_dcacheRW_rdata[9:0] : info_5; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_390 = 4'h6 == select_r ? io_dcacheRW_rdata[9:0] : info_6; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_391 = 4'h7 == select_r ? io_dcacheRW_rdata[9:0] : info_7; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_392 = 4'h8 == select_r ? io_dcacheRW_rdata[9:0] : info_8; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_393 = 4'h9 == select_r ? io_dcacheRW_rdata[9:0] : info_9; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_394 = 4'ha == select_r ? io_dcacheRW_rdata[9:0] : info_10; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_395 = 4'hb == select_r ? io_dcacheRW_rdata[9:0] : info_11; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_396 = 4'hc == select_r ? io_dcacheRW_rdata[9:0] : info_12; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_397 = 4'hd == select_r ? io_dcacheRW_rdata[9:0] : info_13; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_398 = 4'he == select_r ? io_dcacheRW_rdata[9:0] : info_14; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire [9:0] _GEN_399 = 4'hf == select_r ? io_dcacheRW_rdata[9:0] : info_15; // @[tlb.scala 226:40 tlb.scala 226:40 tlb.scala 41:26]
  wire  _GEN_401 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     | _GEN_151; // @[tlb.scala 213:117 tlb.scala 216:40]
  wire [51:0] _GEN_402 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_0 : _GEN_304; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_403 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_1 : _GEN_305; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_404 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_2 : _GEN_306; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_405 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_3 : _GEN_307; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_406 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_4 : _GEN_308; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_407 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_5 : _GEN_309; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_408 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_6 : _GEN_310; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_409 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_7 : _GEN_311; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_410 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_8 : _GEN_312; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_411 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_9 : _GEN_313; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_412 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_10 : _GEN_314; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_413 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_11 : _GEN_315; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_414 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_12 : _GEN_316; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_415 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_13 : _GEN_317; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_416 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_14 : _GEN_318; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire [51:0] _GEN_417 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_15 : _GEN_319; // @[tlb.scala 213:117 tlb.scala 39:26]
  wire  _GEN_418 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_130 : _GEN_320; // @[tlb.scala 213:117]
  wire  _GEN_419 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_131 : _GEN_321; // @[tlb.scala 213:117]
  wire  _GEN_420 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_132 : _GEN_322; // @[tlb.scala 213:117]
  wire  _GEN_421 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_133 : _GEN_323; // @[tlb.scala 213:117]
  wire  _GEN_422 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_134 : _GEN_324; // @[tlb.scala 213:117]
  wire  _GEN_423 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_135 : _GEN_325; // @[tlb.scala 213:117]
  wire  _GEN_424 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_136 : _GEN_326; // @[tlb.scala 213:117]
  wire  _GEN_425 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_137 : _GEN_327; // @[tlb.scala 213:117]
  wire  _GEN_426 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_138 : _GEN_328; // @[tlb.scala 213:117]
  wire  _GEN_427 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_139 : _GEN_329; // @[tlb.scala 213:117]
  wire  _GEN_428 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_140 : _GEN_330; // @[tlb.scala 213:117]
  wire  _GEN_429 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_141 : _GEN_331; // @[tlb.scala 213:117]
  wire  _GEN_430 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_142 : _GEN_332; // @[tlb.scala 213:117]
  wire  _GEN_431 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_143 : _GEN_333; // @[tlb.scala 213:117]
  wire  _GEN_432 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_144 : _GEN_334; // @[tlb.scala 213:117]
  wire  _GEN_433 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_145 : _GEN_335; // @[tlb.scala 213:117]
  wire [19:0] _GEN_434 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_0 : _GEN_336; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_435 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_1 : _GEN_337; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_436 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_2 : _GEN_338; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_437 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_3 : _GEN_339; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_438 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_4 : _GEN_340; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_439 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_5 : _GEN_341; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_440 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_6 : _GEN_342; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_441 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_7 : _GEN_343; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_442 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_8 : _GEN_344; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_443 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_9 : _GEN_345; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_444 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_10 : _GEN_346; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_445 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_11 : _GEN_347; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_446 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_12 : _GEN_348; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_447 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_13 : _GEN_349; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_448 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_14 : _GEN_350; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [19:0] _GEN_449 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_15 : _GEN_351; // @[tlb.scala 213:117 tlb.scala 40:26]
  wire [31:0] _GEN_450 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_0 : _GEN_352; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_451 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_1 : _GEN_353; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_452 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_2 : _GEN_354; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_453 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_3 : _GEN_355; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_454 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_4 : _GEN_356; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_455 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_5 : _GEN_357; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_456 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_6 : _GEN_358; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_457 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_7 : _GEN_359; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_458 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_8 : _GEN_360; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_459 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_9 : _GEN_361; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_460 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_10 : _GEN_362; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_461 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_11 : _GEN_363; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_462 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_12 : _GEN_364; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_463 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_13 : _GEN_365; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_464 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_14 : _GEN_366; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [31:0] _GEN_465 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_15 : _GEN_367; // @[tlb.scala 213:117 tlb.scala 42:30]
  wire [1:0] _GEN_466 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_0 : _GEN_368; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_467 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_1 : _GEN_369; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_468 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_2 : _GEN_370; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_469 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_3 : _GEN_371; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_470 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_4 : _GEN_372; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_471 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_5 : _GEN_373; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_472 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_6 : _GEN_374; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_473 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_7 : _GEN_375; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_474 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_8 : _GEN_376; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_475 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_9 : _GEN_377; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_476 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_10 : _GEN_378; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_477 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_11 : _GEN_379; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_478 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_12 : _GEN_380; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_479 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_13 : _GEN_381; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_480 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_14 : _GEN_382; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [1:0] _GEN_481 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_15 : _GEN_383; // @[tlb.scala 213:117 tlb.scala 43:30]
  wire [9:0] _GEN_482 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_0 : _GEN_384; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_483 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_1 : _GEN_385; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_484 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_2 : _GEN_386; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_485 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_3 : _GEN_387; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_486 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_4 : _GEN_388; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_487 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_5 : _GEN_389; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_488 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_6 : _GEN_390; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_489 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_7 : _GEN_391; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_490 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_8 : _GEN_392; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_491 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_9 : _GEN_393; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_492 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_10 : _GEN_394; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_493 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_11 : _GEN_395; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_494 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_12 : _GEN_396; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_495 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_13 : _GEN_397; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_496 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_14 : _GEN_398; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire [9:0] _GEN_497 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_15 : _GEN_399; // @[tlb.scala 213:117 tlb.scala 41:26]
  wire  _GEN_499 = _T_112 | _GEN_401; // @[tlb.scala 209:99 tlb.scala 212:40]
  wire [51:0] _GEN_500 = _T_112 ? tag_0 : _GEN_402; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_501 = _T_112 ? tag_1 : _GEN_403; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_502 = _T_112 ? tag_2 : _GEN_404; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_503 = _T_112 ? tag_3 : _GEN_405; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_504 = _T_112 ? tag_4 : _GEN_406; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_505 = _T_112 ? tag_5 : _GEN_407; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_506 = _T_112 ? tag_6 : _GEN_408; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_507 = _T_112 ? tag_7 : _GEN_409; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_508 = _T_112 ? tag_8 : _GEN_410; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_509 = _T_112 ? tag_9 : _GEN_411; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_510 = _T_112 ? tag_10 : _GEN_412; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_511 = _T_112 ? tag_11 : _GEN_413; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_512 = _T_112 ? tag_12 : _GEN_414; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_513 = _T_112 ? tag_13 : _GEN_415; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_514 = _T_112 ? tag_14 : _GEN_416; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire [51:0] _GEN_515 = _T_112 ? tag_15 : _GEN_417; // @[tlb.scala 209:99 tlb.scala 39:26]
  wire  _GEN_516 = _T_112 ? _GEN_130 : _GEN_418; // @[tlb.scala 209:99]
  wire  _GEN_517 = _T_112 ? _GEN_131 : _GEN_419; // @[tlb.scala 209:99]
  wire  _GEN_518 = _T_112 ? _GEN_132 : _GEN_420; // @[tlb.scala 209:99]
  wire  _GEN_519 = _T_112 ? _GEN_133 : _GEN_421; // @[tlb.scala 209:99]
  wire  _GEN_520 = _T_112 ? _GEN_134 : _GEN_422; // @[tlb.scala 209:99]
  wire  _GEN_521 = _T_112 ? _GEN_135 : _GEN_423; // @[tlb.scala 209:99]
  wire  _GEN_522 = _T_112 ? _GEN_136 : _GEN_424; // @[tlb.scala 209:99]
  wire  _GEN_523 = _T_112 ? _GEN_137 : _GEN_425; // @[tlb.scala 209:99]
  wire  _GEN_524 = _T_112 ? _GEN_138 : _GEN_426; // @[tlb.scala 209:99]
  wire  _GEN_525 = _T_112 ? _GEN_139 : _GEN_427; // @[tlb.scala 209:99]
  wire  _GEN_526 = _T_112 ? _GEN_140 : _GEN_428; // @[tlb.scala 209:99]
  wire  _GEN_527 = _T_112 ? _GEN_141 : _GEN_429; // @[tlb.scala 209:99]
  wire  _GEN_528 = _T_112 ? _GEN_142 : _GEN_430; // @[tlb.scala 209:99]
  wire  _GEN_529 = _T_112 ? _GEN_143 : _GEN_431; // @[tlb.scala 209:99]
  wire  _GEN_530 = _T_112 ? _GEN_144 : _GEN_432; // @[tlb.scala 209:99]
  wire  _GEN_531 = _T_112 ? _GEN_145 : _GEN_433; // @[tlb.scala 209:99]
  wire [19:0] _GEN_532 = _T_112 ? paddr_0 : _GEN_434; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_533 = _T_112 ? paddr_1 : _GEN_435; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_534 = _T_112 ? paddr_2 : _GEN_436; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_535 = _T_112 ? paddr_3 : _GEN_437; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_536 = _T_112 ? paddr_4 : _GEN_438; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_537 = _T_112 ? paddr_5 : _GEN_439; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_538 = _T_112 ? paddr_6 : _GEN_440; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_539 = _T_112 ? paddr_7 : _GEN_441; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_540 = _T_112 ? paddr_8 : _GEN_442; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_541 = _T_112 ? paddr_9 : _GEN_443; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_542 = _T_112 ? paddr_10 : _GEN_444; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_543 = _T_112 ? paddr_11 : _GEN_445; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_544 = _T_112 ? paddr_12 : _GEN_446; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_545 = _T_112 ? paddr_13 : _GEN_447; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_546 = _T_112 ? paddr_14 : _GEN_448; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [19:0] _GEN_547 = _T_112 ? paddr_15 : _GEN_449; // @[tlb.scala 209:99 tlb.scala 40:26]
  wire [31:0] _GEN_548 = _T_112 ? pte_addr_0 : _GEN_450; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_549 = _T_112 ? pte_addr_1 : _GEN_451; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_550 = _T_112 ? pte_addr_2 : _GEN_452; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_551 = _T_112 ? pte_addr_3 : _GEN_453; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_552 = _T_112 ? pte_addr_4 : _GEN_454; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_553 = _T_112 ? pte_addr_5 : _GEN_455; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_554 = _T_112 ? pte_addr_6 : _GEN_456; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_555 = _T_112 ? pte_addr_7 : _GEN_457; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_556 = _T_112 ? pte_addr_8 : _GEN_458; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_557 = _T_112 ? pte_addr_9 : _GEN_459; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_558 = _T_112 ? pte_addr_10 : _GEN_460; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_559 = _T_112 ? pte_addr_11 : _GEN_461; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_560 = _T_112 ? pte_addr_12 : _GEN_462; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_561 = _T_112 ? pte_addr_13 : _GEN_463; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_562 = _T_112 ? pte_addr_14 : _GEN_464; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [31:0] _GEN_563 = _T_112 ? pte_addr_15 : _GEN_465; // @[tlb.scala 209:99 tlb.scala 42:30]
  wire [1:0] _GEN_564 = _T_112 ? pte_level_0 : _GEN_466; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_565 = _T_112 ? pte_level_1 : _GEN_467; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_566 = _T_112 ? pte_level_2 : _GEN_468; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_567 = _T_112 ? pte_level_3 : _GEN_469; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_568 = _T_112 ? pte_level_4 : _GEN_470; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_569 = _T_112 ? pte_level_5 : _GEN_471; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_570 = _T_112 ? pte_level_6 : _GEN_472; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_571 = _T_112 ? pte_level_7 : _GEN_473; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_572 = _T_112 ? pte_level_8 : _GEN_474; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_573 = _T_112 ? pte_level_9 : _GEN_475; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_574 = _T_112 ? pte_level_10 : _GEN_476; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_575 = _T_112 ? pte_level_11 : _GEN_477; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_576 = _T_112 ? pte_level_12 : _GEN_478; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_577 = _T_112 ? pte_level_13 : _GEN_479; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_578 = _T_112 ? pte_level_14 : _GEN_480; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [1:0] _GEN_579 = _T_112 ? pte_level_15 : _GEN_481; // @[tlb.scala 209:99 tlb.scala 43:30]
  wire [9:0] _GEN_580 = _T_112 ? info_0 : _GEN_482; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_581 = _T_112 ? info_1 : _GEN_483; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_582 = _T_112 ? info_2 : _GEN_484; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_583 = _T_112 ? info_3 : _GEN_485; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_584 = _T_112 ? info_4 : _GEN_486; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_585 = _T_112 ? info_5 : _GEN_487; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_586 = _T_112 ? info_6 : _GEN_488; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_587 = _T_112 ? info_7 : _GEN_489; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_588 = _T_112 ? info_8 : _GEN_490; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_589 = _T_112 ? info_9 : _GEN_491; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_590 = _T_112 ? info_10 : _GEN_492; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_591 = _T_112 ? info_11 : _GEN_493; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_592 = _T_112 ? info_12 : _GEN_494; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_593 = _T_112 ? info_13 : _GEN_495; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_594 = _T_112 ? info_14 : _GEN_496; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire [9:0] _GEN_595 = _T_112 ? info_15 : _GEN_497; // @[tlb.scala 209:99 tlb.scala 41:26]
  wire  _GEN_597 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] | _GEN_499; // @[tlb.scala 203:87 tlb.scala 206:40]
  wire [51:0] _GEN_598 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_0 : _GEN_500; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_599 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_1 : _GEN_501; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_600 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_2 : _GEN_502; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_601 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_3 : _GEN_503; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_602 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_4 : _GEN_504; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_603 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_5 : _GEN_505; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_604 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_6 : _GEN_506; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_605 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_7 : _GEN_507; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_606 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_8 : _GEN_508; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_607 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_9 : _GEN_509; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_608 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_10 : _GEN_510; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_609 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_11 : _GEN_511; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_610 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_12 : _GEN_512; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_611 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_13 : _GEN_513; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_612 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_14 : _GEN_514; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire [51:0] _GEN_613 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_15 : _GEN_515; // @[tlb.scala 203:87 tlb.scala 39:26]
  wire  _GEN_614 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_130 : _GEN_516; // @[tlb.scala 203:87]
  wire  _GEN_615 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_131 : _GEN_517; // @[tlb.scala 203:87]
  wire  _GEN_616 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_132 : _GEN_518; // @[tlb.scala 203:87]
  wire  _GEN_617 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_133 : _GEN_519; // @[tlb.scala 203:87]
  wire  _GEN_618 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_134 : _GEN_520; // @[tlb.scala 203:87]
  wire  _GEN_619 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_135 : _GEN_521; // @[tlb.scala 203:87]
  wire  _GEN_620 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_136 : _GEN_522; // @[tlb.scala 203:87]
  wire  _GEN_621 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_137 : _GEN_523; // @[tlb.scala 203:87]
  wire  _GEN_622 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_138 : _GEN_524; // @[tlb.scala 203:87]
  wire  _GEN_623 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_139 : _GEN_525; // @[tlb.scala 203:87]
  wire  _GEN_624 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_140 : _GEN_526; // @[tlb.scala 203:87]
  wire  _GEN_625 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_141 : _GEN_527; // @[tlb.scala 203:87]
  wire  _GEN_626 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_142 : _GEN_528; // @[tlb.scala 203:87]
  wire  _GEN_627 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_143 : _GEN_529; // @[tlb.scala 203:87]
  wire  _GEN_628 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_144 : _GEN_530; // @[tlb.scala 203:87]
  wire  _GEN_629 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_145 : _GEN_531; // @[tlb.scala 203:87]
  wire [19:0] _GEN_630 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_0 : _GEN_532; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_631 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_1 : _GEN_533; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_632 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_2 : _GEN_534; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_633 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_3 : _GEN_535; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_634 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_4 : _GEN_536; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_635 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_5 : _GEN_537; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_636 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_6 : _GEN_538; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_637 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_7 : _GEN_539; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_638 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_8 : _GEN_540; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_639 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_9 : _GEN_541; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_640 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_10 : _GEN_542; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_641 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_11 : _GEN_543; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_642 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_12 : _GEN_544; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_643 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_13 : _GEN_545; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_644 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_14 : _GEN_546; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [19:0] _GEN_645 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_15 : _GEN_547; // @[tlb.scala 203:87 tlb.scala 40:26]
  wire [31:0] _GEN_646 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_0 : _GEN_548; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_647 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_1 : _GEN_549; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_648 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_2 : _GEN_550; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_649 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_3 : _GEN_551; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_650 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_4 : _GEN_552; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_651 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_5 : _GEN_553; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_652 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_6 : _GEN_554; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_653 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_7 : _GEN_555; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_654 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_8 : _GEN_556; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_655 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_9 : _GEN_557; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_656 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_10 : _GEN_558; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_657 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_11 : _GEN_559; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_658 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_12 : _GEN_560; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_659 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_13 : _GEN_561; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_660 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_14 : _GEN_562; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [31:0] _GEN_661 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_15 : _GEN_563; // @[tlb.scala 203:87 tlb.scala 42:30]
  wire [1:0] _GEN_662 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_0 : _GEN_564; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_663 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_1 : _GEN_565; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_664 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_2 : _GEN_566; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_665 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_3 : _GEN_567; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_666 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_4 : _GEN_568; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_667 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_5 : _GEN_569; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_668 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_6 : _GEN_570; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_669 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_7 : _GEN_571; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_670 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_8 : _GEN_572; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_671 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_9 : _GEN_573; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_672 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_10 : _GEN_574; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_673 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_11 : _GEN_575; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_674 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_12 : _GEN_576; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_675 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_13 : _GEN_577; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_676 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_14 : _GEN_578; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [1:0] _GEN_677 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_15 : _GEN_579; // @[tlb.scala 203:87 tlb.scala 43:30]
  wire [9:0] _GEN_678 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_0 : _GEN_580; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_679 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_1 : _GEN_581; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_680 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_2 : _GEN_582; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_681 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_3 : _GEN_583; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_682 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_4 : _GEN_584; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_683 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_5 : _GEN_585; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_684 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_6 : _GEN_586; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_685 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_7 : _GEN_587; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_686 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_8 : _GEN_588; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_687 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_9 : _GEN_589; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_688 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_10 : _GEN_590; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_689 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_11 : _GEN_591; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_690 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_12 : _GEN_592; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_691 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_13 : _GEN_593; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_692 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_14 : _GEN_594; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire [9:0] _GEN_693 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_15 : _GEN_595; // @[tlb.scala 203:87 tlb.scala 41:26]
  wire  _GEN_695 = _T_87 | _GEN_597; // @[tlb.scala 199:193 tlb.scala 202:40]
  wire [51:0] _GEN_696 = _T_87 ? tag_0 : _GEN_598; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_697 = _T_87 ? tag_1 : _GEN_599; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_698 = _T_87 ? tag_2 : _GEN_600; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_699 = _T_87 ? tag_3 : _GEN_601; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_700 = _T_87 ? tag_4 : _GEN_602; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_701 = _T_87 ? tag_5 : _GEN_603; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_702 = _T_87 ? tag_6 : _GEN_604; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_703 = _T_87 ? tag_7 : _GEN_605; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_704 = _T_87 ? tag_8 : _GEN_606; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_705 = _T_87 ? tag_9 : _GEN_607; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_706 = _T_87 ? tag_10 : _GEN_608; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_707 = _T_87 ? tag_11 : _GEN_609; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_708 = _T_87 ? tag_12 : _GEN_610; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_709 = _T_87 ? tag_13 : _GEN_611; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_710 = _T_87 ? tag_14 : _GEN_612; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire [51:0] _GEN_711 = _T_87 ? tag_15 : _GEN_613; // @[tlb.scala 199:193 tlb.scala 39:26]
  wire  _GEN_712 = _T_87 ? _GEN_130 : _GEN_614; // @[tlb.scala 199:193]
  wire  _GEN_713 = _T_87 ? _GEN_131 : _GEN_615; // @[tlb.scala 199:193]
  wire  _GEN_714 = _T_87 ? _GEN_132 : _GEN_616; // @[tlb.scala 199:193]
  wire  _GEN_715 = _T_87 ? _GEN_133 : _GEN_617; // @[tlb.scala 199:193]
  wire  _GEN_716 = _T_87 ? _GEN_134 : _GEN_618; // @[tlb.scala 199:193]
  wire  _GEN_717 = _T_87 ? _GEN_135 : _GEN_619; // @[tlb.scala 199:193]
  wire  _GEN_718 = _T_87 ? _GEN_136 : _GEN_620; // @[tlb.scala 199:193]
  wire  _GEN_719 = _T_87 ? _GEN_137 : _GEN_621; // @[tlb.scala 199:193]
  wire  _GEN_720 = _T_87 ? _GEN_138 : _GEN_622; // @[tlb.scala 199:193]
  wire  _GEN_721 = _T_87 ? _GEN_139 : _GEN_623; // @[tlb.scala 199:193]
  wire  _GEN_722 = _T_87 ? _GEN_140 : _GEN_624; // @[tlb.scala 199:193]
  wire  _GEN_723 = _T_87 ? _GEN_141 : _GEN_625; // @[tlb.scala 199:193]
  wire  _GEN_724 = _T_87 ? _GEN_142 : _GEN_626; // @[tlb.scala 199:193]
  wire  _GEN_725 = _T_87 ? _GEN_143 : _GEN_627; // @[tlb.scala 199:193]
  wire  _GEN_726 = _T_87 ? _GEN_144 : _GEN_628; // @[tlb.scala 199:193]
  wire  _GEN_727 = _T_87 ? _GEN_145 : _GEN_629; // @[tlb.scala 199:193]
  wire [19:0] _GEN_728 = _T_87 ? paddr_0 : _GEN_630; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_729 = _T_87 ? paddr_1 : _GEN_631; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_730 = _T_87 ? paddr_2 : _GEN_632; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_731 = _T_87 ? paddr_3 : _GEN_633; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_732 = _T_87 ? paddr_4 : _GEN_634; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_733 = _T_87 ? paddr_5 : _GEN_635; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_734 = _T_87 ? paddr_6 : _GEN_636; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_735 = _T_87 ? paddr_7 : _GEN_637; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_736 = _T_87 ? paddr_8 : _GEN_638; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_737 = _T_87 ? paddr_9 : _GEN_639; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_738 = _T_87 ? paddr_10 : _GEN_640; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_739 = _T_87 ? paddr_11 : _GEN_641; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_740 = _T_87 ? paddr_12 : _GEN_642; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_741 = _T_87 ? paddr_13 : _GEN_643; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_742 = _T_87 ? paddr_14 : _GEN_644; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [19:0] _GEN_743 = _T_87 ? paddr_15 : _GEN_645; // @[tlb.scala 199:193 tlb.scala 40:26]
  wire [31:0] _GEN_744 = _T_87 ? pte_addr_0 : _GEN_646; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_745 = _T_87 ? pte_addr_1 : _GEN_647; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_746 = _T_87 ? pte_addr_2 : _GEN_648; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_747 = _T_87 ? pte_addr_3 : _GEN_649; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_748 = _T_87 ? pte_addr_4 : _GEN_650; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_749 = _T_87 ? pte_addr_5 : _GEN_651; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_750 = _T_87 ? pte_addr_6 : _GEN_652; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_751 = _T_87 ? pte_addr_7 : _GEN_653; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_752 = _T_87 ? pte_addr_8 : _GEN_654; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_753 = _T_87 ? pte_addr_9 : _GEN_655; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_754 = _T_87 ? pte_addr_10 : _GEN_656; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_755 = _T_87 ? pte_addr_11 : _GEN_657; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_756 = _T_87 ? pte_addr_12 : _GEN_658; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_757 = _T_87 ? pte_addr_13 : _GEN_659; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_758 = _T_87 ? pte_addr_14 : _GEN_660; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [31:0] _GEN_759 = _T_87 ? pte_addr_15 : _GEN_661; // @[tlb.scala 199:193 tlb.scala 42:30]
  wire [1:0] _GEN_760 = _T_87 ? pte_level_0 : _GEN_662; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_761 = _T_87 ? pte_level_1 : _GEN_663; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_762 = _T_87 ? pte_level_2 : _GEN_664; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_763 = _T_87 ? pte_level_3 : _GEN_665; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_764 = _T_87 ? pte_level_4 : _GEN_666; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_765 = _T_87 ? pte_level_5 : _GEN_667; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_766 = _T_87 ? pte_level_6 : _GEN_668; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_767 = _T_87 ? pte_level_7 : _GEN_669; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_768 = _T_87 ? pte_level_8 : _GEN_670; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_769 = _T_87 ? pte_level_9 : _GEN_671; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_770 = _T_87 ? pte_level_10 : _GEN_672; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_771 = _T_87 ? pte_level_11 : _GEN_673; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_772 = _T_87 ? pte_level_12 : _GEN_674; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_773 = _T_87 ? pte_level_13 : _GEN_675; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_774 = _T_87 ? pte_level_14 : _GEN_676; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [1:0] _GEN_775 = _T_87 ? pte_level_15 : _GEN_677; // @[tlb.scala 199:193 tlb.scala 43:30]
  wire [9:0] _GEN_776 = _T_87 ? info_0 : _GEN_678; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_777 = _T_87 ? info_1 : _GEN_679; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_778 = _T_87 ? info_2 : _GEN_680; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_779 = _T_87 ? info_3 : _GEN_681; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_780 = _T_87 ? info_4 : _GEN_682; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_781 = _T_87 ? info_5 : _GEN_683; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_782 = _T_87 ? info_6 : _GEN_684; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_783 = _T_87 ? info_7 : _GEN_685; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_784 = _T_87 ? info_8 : _GEN_686; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_785 = _T_87 ? info_9 : _GEN_687; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_786 = _T_87 ? info_10 : _GEN_688; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_787 = _T_87 ? info_11 : _GEN_689; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_788 = _T_87 ? info_12 : _GEN_690; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_789 = _T_87 ? info_13 : _GEN_691; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_790 = _T_87 ? info_14 : _GEN_692; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [9:0] _GEN_791 = _T_87 ? info_15 : _GEN_693; // @[tlb.scala 199:193 tlb.scala 41:26]
  wire [1:0] _GEN_792 = _T_73 == 64'h1 ? _GEN_300 : 2'h0; // @[tlb.scala 191:76]
  wire  _GEN_793 = _T_73 == 64'h1 ? _GEN_301 : _GEN_695; // @[tlb.scala 191:76]
  wire [55:0] _GEN_794 = _T_73 == 64'h1 ? _GEN_302 : {{24'd0}, pte_addr_r}; // @[tlb.scala 191:76 tlb.scala 47:30]
  wire [4:0] _GEN_795 = _T_73 == 64'h1 ? _GEN_303 : _GEN_297; // @[tlb.scala 191:76]
  wire [51:0] _GEN_796 = _T_73 == 64'h1 ? tag_0 : _GEN_696; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_797 = _T_73 == 64'h1 ? tag_1 : _GEN_697; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_798 = _T_73 == 64'h1 ? tag_2 : _GEN_698; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_799 = _T_73 == 64'h1 ? tag_3 : _GEN_699; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_800 = _T_73 == 64'h1 ? tag_4 : _GEN_700; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_801 = _T_73 == 64'h1 ? tag_5 : _GEN_701; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_802 = _T_73 == 64'h1 ? tag_6 : _GEN_702; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_803 = _T_73 == 64'h1 ? tag_7 : _GEN_703; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_804 = _T_73 == 64'h1 ? tag_8 : _GEN_704; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_805 = _T_73 == 64'h1 ? tag_9 : _GEN_705; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_806 = _T_73 == 64'h1 ? tag_10 : _GEN_706; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_807 = _T_73 == 64'h1 ? tag_11 : _GEN_707; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_808 = _T_73 == 64'h1 ? tag_12 : _GEN_708; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_809 = _T_73 == 64'h1 ? tag_13 : _GEN_709; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_810 = _T_73 == 64'h1 ? tag_14 : _GEN_710; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire [51:0] _GEN_811 = _T_73 == 64'h1 ? tag_15 : _GEN_711; // @[tlb.scala 191:76 tlb.scala 39:26]
  wire  _GEN_812 = _T_73 == 64'h1 ? _GEN_130 : _GEN_712; // @[tlb.scala 191:76]
  wire  _GEN_813 = _T_73 == 64'h1 ? _GEN_131 : _GEN_713; // @[tlb.scala 191:76]
  wire  _GEN_814 = _T_73 == 64'h1 ? _GEN_132 : _GEN_714; // @[tlb.scala 191:76]
  wire  _GEN_815 = _T_73 == 64'h1 ? _GEN_133 : _GEN_715; // @[tlb.scala 191:76]
  wire  _GEN_816 = _T_73 == 64'h1 ? _GEN_134 : _GEN_716; // @[tlb.scala 191:76]
  wire  _GEN_817 = _T_73 == 64'h1 ? _GEN_135 : _GEN_717; // @[tlb.scala 191:76]
  wire  _GEN_818 = _T_73 == 64'h1 ? _GEN_136 : _GEN_718; // @[tlb.scala 191:76]
  wire  _GEN_819 = _T_73 == 64'h1 ? _GEN_137 : _GEN_719; // @[tlb.scala 191:76]
  wire  _GEN_820 = _T_73 == 64'h1 ? _GEN_138 : _GEN_720; // @[tlb.scala 191:76]
  wire  _GEN_821 = _T_73 == 64'h1 ? _GEN_139 : _GEN_721; // @[tlb.scala 191:76]
  wire  _GEN_822 = _T_73 == 64'h1 ? _GEN_140 : _GEN_722; // @[tlb.scala 191:76]
  wire  _GEN_823 = _T_73 == 64'h1 ? _GEN_141 : _GEN_723; // @[tlb.scala 191:76]
  wire  _GEN_824 = _T_73 == 64'h1 ? _GEN_142 : _GEN_724; // @[tlb.scala 191:76]
  wire  _GEN_825 = _T_73 == 64'h1 ? _GEN_143 : _GEN_725; // @[tlb.scala 191:76]
  wire  _GEN_826 = _T_73 == 64'h1 ? _GEN_144 : _GEN_726; // @[tlb.scala 191:76]
  wire  _GEN_827 = _T_73 == 64'h1 ? _GEN_145 : _GEN_727; // @[tlb.scala 191:76]
  wire [19:0] _GEN_828 = _T_73 == 64'h1 ? paddr_0 : _GEN_728; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_829 = _T_73 == 64'h1 ? paddr_1 : _GEN_729; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_830 = _T_73 == 64'h1 ? paddr_2 : _GEN_730; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_831 = _T_73 == 64'h1 ? paddr_3 : _GEN_731; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_832 = _T_73 == 64'h1 ? paddr_4 : _GEN_732; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_833 = _T_73 == 64'h1 ? paddr_5 : _GEN_733; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_834 = _T_73 == 64'h1 ? paddr_6 : _GEN_734; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_835 = _T_73 == 64'h1 ? paddr_7 : _GEN_735; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_836 = _T_73 == 64'h1 ? paddr_8 : _GEN_736; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_837 = _T_73 == 64'h1 ? paddr_9 : _GEN_737; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_838 = _T_73 == 64'h1 ? paddr_10 : _GEN_738; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_839 = _T_73 == 64'h1 ? paddr_11 : _GEN_739; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_840 = _T_73 == 64'h1 ? paddr_12 : _GEN_740; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_841 = _T_73 == 64'h1 ? paddr_13 : _GEN_741; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_842 = _T_73 == 64'h1 ? paddr_14 : _GEN_742; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [19:0] _GEN_843 = _T_73 == 64'h1 ? paddr_15 : _GEN_743; // @[tlb.scala 191:76 tlb.scala 40:26]
  wire [31:0] _GEN_844 = _T_73 == 64'h1 ? pte_addr_0 : _GEN_744; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_845 = _T_73 == 64'h1 ? pte_addr_1 : _GEN_745; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_846 = _T_73 == 64'h1 ? pte_addr_2 : _GEN_746; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_847 = _T_73 == 64'h1 ? pte_addr_3 : _GEN_747; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_848 = _T_73 == 64'h1 ? pte_addr_4 : _GEN_748; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_849 = _T_73 == 64'h1 ? pte_addr_5 : _GEN_749; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_850 = _T_73 == 64'h1 ? pte_addr_6 : _GEN_750; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_851 = _T_73 == 64'h1 ? pte_addr_7 : _GEN_751; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_852 = _T_73 == 64'h1 ? pte_addr_8 : _GEN_752; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_853 = _T_73 == 64'h1 ? pte_addr_9 : _GEN_753; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_854 = _T_73 == 64'h1 ? pte_addr_10 : _GEN_754; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_855 = _T_73 == 64'h1 ? pte_addr_11 : _GEN_755; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_856 = _T_73 == 64'h1 ? pte_addr_12 : _GEN_756; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_857 = _T_73 == 64'h1 ? pte_addr_13 : _GEN_757; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_858 = _T_73 == 64'h1 ? pte_addr_14 : _GEN_758; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [31:0] _GEN_859 = _T_73 == 64'h1 ? pte_addr_15 : _GEN_759; // @[tlb.scala 191:76 tlb.scala 42:30]
  wire [1:0] _GEN_860 = _T_73 == 64'h1 ? pte_level_0 : _GEN_760; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_861 = _T_73 == 64'h1 ? pte_level_1 : _GEN_761; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_862 = _T_73 == 64'h1 ? pte_level_2 : _GEN_762; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_863 = _T_73 == 64'h1 ? pte_level_3 : _GEN_763; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_864 = _T_73 == 64'h1 ? pte_level_4 : _GEN_764; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_865 = _T_73 == 64'h1 ? pte_level_5 : _GEN_765; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_866 = _T_73 == 64'h1 ? pte_level_6 : _GEN_766; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_867 = _T_73 == 64'h1 ? pte_level_7 : _GEN_767; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_868 = _T_73 == 64'h1 ? pte_level_8 : _GEN_768; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_869 = _T_73 == 64'h1 ? pte_level_9 : _GEN_769; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_870 = _T_73 == 64'h1 ? pte_level_10 : _GEN_770; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_871 = _T_73 == 64'h1 ? pte_level_11 : _GEN_771; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_872 = _T_73 == 64'h1 ? pte_level_12 : _GEN_772; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_873 = _T_73 == 64'h1 ? pte_level_13 : _GEN_773; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_874 = _T_73 == 64'h1 ? pte_level_14 : _GEN_774; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [1:0] _GEN_875 = _T_73 == 64'h1 ? pte_level_15 : _GEN_775; // @[tlb.scala 191:76 tlb.scala 43:30]
  wire [9:0] _GEN_876 = _T_73 == 64'h1 ? info_0 : _GEN_776; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_877 = _T_73 == 64'h1 ? info_1 : _GEN_777; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_878 = _T_73 == 64'h1 ? info_2 : _GEN_778; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_879 = _T_73 == 64'h1 ? info_3 : _GEN_779; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_880 = _T_73 == 64'h1 ? info_4 : _GEN_780; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_881 = _T_73 == 64'h1 ? info_5 : _GEN_781; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_882 = _T_73 == 64'h1 ? info_6 : _GEN_782; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_883 = _T_73 == 64'h1 ? info_7 : _GEN_783; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_884 = _T_73 == 64'h1 ? info_8 : _GEN_784; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_885 = _T_73 == 64'h1 ? info_9 : _GEN_785; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_886 = _T_73 == 64'h1 ? info_10 : _GEN_786; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_887 = _T_73 == 64'h1 ? info_11 : _GEN_787; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_888 = _T_73 == 64'h1 ? info_12 : _GEN_788; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_889 = _T_73 == 64'h1 ? info_13 : _GEN_789; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_890 = _T_73 == 64'h1 ? info_14 : _GEN_790; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [9:0] _GEN_891 = _T_73 == 64'h1 ? info_15 : _GEN_791; // @[tlb.scala 191:76 tlb.scala 41:26]
  wire [1:0] _GEN_892 = io_dcacheRW_rvalid ? _GEN_792 : state; // @[tlb.scala 190:41 tlb.scala 84:24]
  wire  _GEN_893 = io_dcacheRW_rvalid ? _GEN_793 : _GEN_151; // @[tlb.scala 190:41]
  wire [55:0] _GEN_894 = io_dcacheRW_rvalid ? _GEN_794 : {{24'd0}, pte_addr_r}; // @[tlb.scala 190:41 tlb.scala 47:30]
  wire [4:0] _GEN_895 = io_dcacheRW_rvalid ? _GEN_795 : _GEN_297; // @[tlb.scala 190:41]
  wire [51:0] _GEN_896 = io_dcacheRW_rvalid ? _GEN_796 : tag_0; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_897 = io_dcacheRW_rvalid ? _GEN_797 : tag_1; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_898 = io_dcacheRW_rvalid ? _GEN_798 : tag_2; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_899 = io_dcacheRW_rvalid ? _GEN_799 : tag_3; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_900 = io_dcacheRW_rvalid ? _GEN_800 : tag_4; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_901 = io_dcacheRW_rvalid ? _GEN_801 : tag_5; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_902 = io_dcacheRW_rvalid ? _GEN_802 : tag_6; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_903 = io_dcacheRW_rvalid ? _GEN_803 : tag_7; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_904 = io_dcacheRW_rvalid ? _GEN_804 : tag_8; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_905 = io_dcacheRW_rvalid ? _GEN_805 : tag_9; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_906 = io_dcacheRW_rvalid ? _GEN_806 : tag_10; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_907 = io_dcacheRW_rvalid ? _GEN_807 : tag_11; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_908 = io_dcacheRW_rvalid ? _GEN_808 : tag_12; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_909 = io_dcacheRW_rvalid ? _GEN_809 : tag_13; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_910 = io_dcacheRW_rvalid ? _GEN_810 : tag_14; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire [51:0] _GEN_911 = io_dcacheRW_rvalid ? _GEN_811 : tag_15; // @[tlb.scala 190:41 tlb.scala 39:26]
  wire  _GEN_912 = io_dcacheRW_rvalid ? _GEN_812 : _GEN_130; // @[tlb.scala 190:41]
  wire  _GEN_913 = io_dcacheRW_rvalid ? _GEN_813 : _GEN_131; // @[tlb.scala 190:41]
  wire  _GEN_914 = io_dcacheRW_rvalid ? _GEN_814 : _GEN_132; // @[tlb.scala 190:41]
  wire  _GEN_915 = io_dcacheRW_rvalid ? _GEN_815 : _GEN_133; // @[tlb.scala 190:41]
  wire  _GEN_916 = io_dcacheRW_rvalid ? _GEN_816 : _GEN_134; // @[tlb.scala 190:41]
  wire  _GEN_917 = io_dcacheRW_rvalid ? _GEN_817 : _GEN_135; // @[tlb.scala 190:41]
  wire  _GEN_918 = io_dcacheRW_rvalid ? _GEN_818 : _GEN_136; // @[tlb.scala 190:41]
  wire  _GEN_919 = io_dcacheRW_rvalid ? _GEN_819 : _GEN_137; // @[tlb.scala 190:41]
  wire  _GEN_920 = io_dcacheRW_rvalid ? _GEN_820 : _GEN_138; // @[tlb.scala 190:41]
  wire  _GEN_921 = io_dcacheRW_rvalid ? _GEN_821 : _GEN_139; // @[tlb.scala 190:41]
  wire  _GEN_922 = io_dcacheRW_rvalid ? _GEN_822 : _GEN_140; // @[tlb.scala 190:41]
  wire  _GEN_923 = io_dcacheRW_rvalid ? _GEN_823 : _GEN_141; // @[tlb.scala 190:41]
  wire  _GEN_924 = io_dcacheRW_rvalid ? _GEN_824 : _GEN_142; // @[tlb.scala 190:41]
  wire  _GEN_925 = io_dcacheRW_rvalid ? _GEN_825 : _GEN_143; // @[tlb.scala 190:41]
  wire  _GEN_926 = io_dcacheRW_rvalid ? _GEN_826 : _GEN_144; // @[tlb.scala 190:41]
  wire  _GEN_927 = io_dcacheRW_rvalid ? _GEN_827 : _GEN_145; // @[tlb.scala 190:41]
  wire [19:0] _GEN_928 = io_dcacheRW_rvalid ? _GEN_828 : paddr_0; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_929 = io_dcacheRW_rvalid ? _GEN_829 : paddr_1; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_930 = io_dcacheRW_rvalid ? _GEN_830 : paddr_2; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_931 = io_dcacheRW_rvalid ? _GEN_831 : paddr_3; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_932 = io_dcacheRW_rvalid ? _GEN_832 : paddr_4; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_933 = io_dcacheRW_rvalid ? _GEN_833 : paddr_5; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_934 = io_dcacheRW_rvalid ? _GEN_834 : paddr_6; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_935 = io_dcacheRW_rvalid ? _GEN_835 : paddr_7; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_936 = io_dcacheRW_rvalid ? _GEN_836 : paddr_8; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_937 = io_dcacheRW_rvalid ? _GEN_837 : paddr_9; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_938 = io_dcacheRW_rvalid ? _GEN_838 : paddr_10; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_939 = io_dcacheRW_rvalid ? _GEN_839 : paddr_11; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_940 = io_dcacheRW_rvalid ? _GEN_840 : paddr_12; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_941 = io_dcacheRW_rvalid ? _GEN_841 : paddr_13; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_942 = io_dcacheRW_rvalid ? _GEN_842 : paddr_14; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [19:0] _GEN_943 = io_dcacheRW_rvalid ? _GEN_843 : paddr_15; // @[tlb.scala 190:41 tlb.scala 40:26]
  wire [31:0] _GEN_944 = io_dcacheRW_rvalid ? _GEN_844 : pte_addr_0; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_945 = io_dcacheRW_rvalid ? _GEN_845 : pte_addr_1; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_946 = io_dcacheRW_rvalid ? _GEN_846 : pte_addr_2; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_947 = io_dcacheRW_rvalid ? _GEN_847 : pte_addr_3; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_948 = io_dcacheRW_rvalid ? _GEN_848 : pte_addr_4; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_949 = io_dcacheRW_rvalid ? _GEN_849 : pte_addr_5; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_950 = io_dcacheRW_rvalid ? _GEN_850 : pte_addr_6; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_951 = io_dcacheRW_rvalid ? _GEN_851 : pte_addr_7; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_952 = io_dcacheRW_rvalid ? _GEN_852 : pte_addr_8; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_953 = io_dcacheRW_rvalid ? _GEN_853 : pte_addr_9; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_954 = io_dcacheRW_rvalid ? _GEN_854 : pte_addr_10; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_955 = io_dcacheRW_rvalid ? _GEN_855 : pte_addr_11; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_956 = io_dcacheRW_rvalid ? _GEN_856 : pte_addr_12; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_957 = io_dcacheRW_rvalid ? _GEN_857 : pte_addr_13; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_958 = io_dcacheRW_rvalid ? _GEN_858 : pte_addr_14; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [31:0] _GEN_959 = io_dcacheRW_rvalid ? _GEN_859 : pte_addr_15; // @[tlb.scala 190:41 tlb.scala 42:30]
  wire [1:0] _GEN_960 = io_dcacheRW_rvalid ? _GEN_860 : pte_level_0; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_961 = io_dcacheRW_rvalid ? _GEN_861 : pte_level_1; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_962 = io_dcacheRW_rvalid ? _GEN_862 : pte_level_2; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_963 = io_dcacheRW_rvalid ? _GEN_863 : pte_level_3; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_964 = io_dcacheRW_rvalid ? _GEN_864 : pte_level_4; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_965 = io_dcacheRW_rvalid ? _GEN_865 : pte_level_5; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_966 = io_dcacheRW_rvalid ? _GEN_866 : pte_level_6; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_967 = io_dcacheRW_rvalid ? _GEN_867 : pte_level_7; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_968 = io_dcacheRW_rvalid ? _GEN_868 : pte_level_8; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_969 = io_dcacheRW_rvalid ? _GEN_869 : pte_level_9; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_970 = io_dcacheRW_rvalid ? _GEN_870 : pte_level_10; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_971 = io_dcacheRW_rvalid ? _GEN_871 : pte_level_11; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_972 = io_dcacheRW_rvalid ? _GEN_872 : pte_level_12; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_973 = io_dcacheRW_rvalid ? _GEN_873 : pte_level_13; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_974 = io_dcacheRW_rvalid ? _GEN_874 : pte_level_14; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [1:0] _GEN_975 = io_dcacheRW_rvalid ? _GEN_875 : pte_level_15; // @[tlb.scala 190:41 tlb.scala 43:30]
  wire [9:0] _GEN_976 = io_dcacheRW_rvalid ? _GEN_876 : info_0; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_977 = io_dcacheRW_rvalid ? _GEN_877 : info_1; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_978 = io_dcacheRW_rvalid ? _GEN_878 : info_2; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_979 = io_dcacheRW_rvalid ? _GEN_879 : info_3; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_980 = io_dcacheRW_rvalid ? _GEN_880 : info_4; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_981 = io_dcacheRW_rvalid ? _GEN_881 : info_5; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_982 = io_dcacheRW_rvalid ? _GEN_882 : info_6; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_983 = io_dcacheRW_rvalid ? _GEN_883 : info_7; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_984 = io_dcacheRW_rvalid ? _GEN_884 : info_8; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_985 = io_dcacheRW_rvalid ? _GEN_885 : info_9; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_986 = io_dcacheRW_rvalid ? _GEN_886 : info_10; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_987 = io_dcacheRW_rvalid ? _GEN_887 : info_11; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_988 = io_dcacheRW_rvalid ? _GEN_888 : info_12; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_989 = io_dcacheRW_rvalid ? _GEN_889 : info_13; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_990 = io_dcacheRW_rvalid ? _GEN_890 : info_14; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [9:0] _GEN_991 = io_dcacheRW_rvalid ? _GEN_891 : info_15; // @[tlb.scala 190:41 tlb.scala 41:26]
  wire [4:0] _GEN_992 = _T_69 ? _GEN_895 : dc_mode_r; // @[Conditional.scala 39:67 tlb.scala 49:30]
  wire [7:0] _GEN_993 = _T_69 ? _GEN_298 : offset; // @[Conditional.scala 39:67 tlb.scala 131:26]
  wire [1:0] _GEN_994 = _T_69 ? _GEN_299 : level; // @[Conditional.scala 39:67 tlb.scala 132:26]
  wire [1:0] _GEN_995 = _T_69 ? _GEN_892 : state; // @[Conditional.scala 39:67 tlb.scala 84:24]
  wire  _GEN_996 = _T_69 ? _GEN_893 : _GEN_151; // @[Conditional.scala 39:67]
  wire [55:0] _GEN_997 = _T_69 ? _GEN_894 : {{24'd0}, pte_addr_r}; // @[Conditional.scala 39:67 tlb.scala 47:30]
  wire [51:0] _GEN_998 = _T_69 ? _GEN_896 : tag_0; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_999 = _T_69 ? _GEN_897 : tag_1; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1000 = _T_69 ? _GEN_898 : tag_2; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1001 = _T_69 ? _GEN_899 : tag_3; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1002 = _T_69 ? _GEN_900 : tag_4; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1003 = _T_69 ? _GEN_901 : tag_5; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1004 = _T_69 ? _GEN_902 : tag_6; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1005 = _T_69 ? _GEN_903 : tag_7; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1006 = _T_69 ? _GEN_904 : tag_8; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1007 = _T_69 ? _GEN_905 : tag_9; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1008 = _T_69 ? _GEN_906 : tag_10; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1009 = _T_69 ? _GEN_907 : tag_11; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1010 = _T_69 ? _GEN_908 : tag_12; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1011 = _T_69 ? _GEN_909 : tag_13; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1012 = _T_69 ? _GEN_910 : tag_14; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire [51:0] _GEN_1013 = _T_69 ? _GEN_911 : tag_15; // @[Conditional.scala 39:67 tlb.scala 39:26]
  wire  _GEN_1014 = _T_69 ? _GEN_912 : _GEN_130; // @[Conditional.scala 39:67]
  wire  _GEN_1015 = _T_69 ? _GEN_913 : _GEN_131; // @[Conditional.scala 39:67]
  wire  _GEN_1016 = _T_69 ? _GEN_914 : _GEN_132; // @[Conditional.scala 39:67]
  wire  _GEN_1017 = _T_69 ? _GEN_915 : _GEN_133; // @[Conditional.scala 39:67]
  wire  _GEN_1018 = _T_69 ? _GEN_916 : _GEN_134; // @[Conditional.scala 39:67]
  wire  _GEN_1019 = _T_69 ? _GEN_917 : _GEN_135; // @[Conditional.scala 39:67]
  wire  _GEN_1020 = _T_69 ? _GEN_918 : _GEN_136; // @[Conditional.scala 39:67]
  wire  _GEN_1021 = _T_69 ? _GEN_919 : _GEN_137; // @[Conditional.scala 39:67]
  wire  _GEN_1022 = _T_69 ? _GEN_920 : _GEN_138; // @[Conditional.scala 39:67]
  wire  _GEN_1023 = _T_69 ? _GEN_921 : _GEN_139; // @[Conditional.scala 39:67]
  wire  _GEN_1024 = _T_69 ? _GEN_922 : _GEN_140; // @[Conditional.scala 39:67]
  wire  _GEN_1025 = _T_69 ? _GEN_923 : _GEN_141; // @[Conditional.scala 39:67]
  wire  _GEN_1026 = _T_69 ? _GEN_924 : _GEN_142; // @[Conditional.scala 39:67]
  wire  _GEN_1027 = _T_69 ? _GEN_925 : _GEN_143; // @[Conditional.scala 39:67]
  wire  _GEN_1028 = _T_69 ? _GEN_926 : _GEN_144; // @[Conditional.scala 39:67]
  wire  _GEN_1029 = _T_69 ? _GEN_927 : _GEN_145; // @[Conditional.scala 39:67]
  wire [19:0] _GEN_1030 = _T_69 ? _GEN_928 : paddr_0; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1031 = _T_69 ? _GEN_929 : paddr_1; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1032 = _T_69 ? _GEN_930 : paddr_2; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1033 = _T_69 ? _GEN_931 : paddr_3; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1034 = _T_69 ? _GEN_932 : paddr_4; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1035 = _T_69 ? _GEN_933 : paddr_5; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1036 = _T_69 ? _GEN_934 : paddr_6; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1037 = _T_69 ? _GEN_935 : paddr_7; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1038 = _T_69 ? _GEN_936 : paddr_8; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1039 = _T_69 ? _GEN_937 : paddr_9; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1040 = _T_69 ? _GEN_938 : paddr_10; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1041 = _T_69 ? _GEN_939 : paddr_11; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1042 = _T_69 ? _GEN_940 : paddr_12; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1043 = _T_69 ? _GEN_941 : paddr_13; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1044 = _T_69 ? _GEN_942 : paddr_14; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [19:0] _GEN_1045 = _T_69 ? _GEN_943 : paddr_15; // @[Conditional.scala 39:67 tlb.scala 40:26]
  wire [31:0] _GEN_1046 = _T_69 ? _GEN_944 : pte_addr_0; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1047 = _T_69 ? _GEN_945 : pte_addr_1; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1048 = _T_69 ? _GEN_946 : pte_addr_2; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1049 = _T_69 ? _GEN_947 : pte_addr_3; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1050 = _T_69 ? _GEN_948 : pte_addr_4; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1051 = _T_69 ? _GEN_949 : pte_addr_5; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1052 = _T_69 ? _GEN_950 : pte_addr_6; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1053 = _T_69 ? _GEN_951 : pte_addr_7; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1054 = _T_69 ? _GEN_952 : pte_addr_8; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1055 = _T_69 ? _GEN_953 : pte_addr_9; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1056 = _T_69 ? _GEN_954 : pte_addr_10; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1057 = _T_69 ? _GEN_955 : pte_addr_11; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1058 = _T_69 ? _GEN_956 : pte_addr_12; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1059 = _T_69 ? _GEN_957 : pte_addr_13; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1060 = _T_69 ? _GEN_958 : pte_addr_14; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [31:0] _GEN_1061 = _T_69 ? _GEN_959 : pte_addr_15; // @[Conditional.scala 39:67 tlb.scala 42:30]
  wire [1:0] _GEN_1062 = _T_69 ? _GEN_960 : pte_level_0; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1063 = _T_69 ? _GEN_961 : pte_level_1; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1064 = _T_69 ? _GEN_962 : pte_level_2; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1065 = _T_69 ? _GEN_963 : pte_level_3; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1066 = _T_69 ? _GEN_964 : pte_level_4; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1067 = _T_69 ? _GEN_965 : pte_level_5; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1068 = _T_69 ? _GEN_966 : pte_level_6; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1069 = _T_69 ? _GEN_967 : pte_level_7; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1070 = _T_69 ? _GEN_968 : pte_level_8; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1071 = _T_69 ? _GEN_969 : pte_level_9; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1072 = _T_69 ? _GEN_970 : pte_level_10; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1073 = _T_69 ? _GEN_971 : pte_level_11; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1074 = _T_69 ? _GEN_972 : pte_level_12; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1075 = _T_69 ? _GEN_973 : pte_level_13; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1076 = _T_69 ? _GEN_974 : pte_level_14; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [1:0] _GEN_1077 = _T_69 ? _GEN_975 : pte_level_15; // @[Conditional.scala 39:67 tlb.scala 43:30]
  wire [9:0] _GEN_1078 = _T_69 ? _GEN_976 : info_0; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1079 = _T_69 ? _GEN_977 : info_1; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1080 = _T_69 ? _GEN_978 : info_2; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1081 = _T_69 ? _GEN_979 : info_3; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1082 = _T_69 ? _GEN_980 : info_4; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1083 = _T_69 ? _GEN_981 : info_5; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1084 = _T_69 ? _GEN_982 : info_6; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1085 = _T_69 ? _GEN_983 : info_7; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1086 = _T_69 ? _GEN_984 : info_8; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1087 = _T_69 ? _GEN_985 : info_9; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1088 = _T_69 ? _GEN_986 : info_10; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1089 = _T_69 ? _GEN_987 : info_11; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1090 = _T_69 ? _GEN_988 : info_12; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1091 = _T_69 ? _GEN_989 : info_13; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1092 = _T_69 ? _GEN_990 : info_14; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [9:0] _GEN_1093 = _T_69 ? _GEN_991 : info_15; // @[Conditional.scala 39:67 tlb.scala 41:26]
  wire [55:0] _GEN_1100 = _T_68 ? {{24'd0}, pte_addr_r} : _GEN_997; // @[Conditional.scala 39:67 tlb.scala 47:30]
  wire [63:0] _GEN_1202 = _T_54 ? _GEN_268 : {{32'd0}, out_paddr_r}; // @[Conditional.scala 40:58 tlb.scala 52:30]
  wire [55:0] _GEN_1205 = _T_54 ? _GEN_271 : _GEN_1100; // @[Conditional.scala 40:58]
  wire [63:0] _GEN_1312 = is_Sv39 | state != 2'h0 ? _GEN_1202 : io_va2pa_vaddr; // @[tlb.scala 135:37 tlb.scala 233:21]
  wire [55:0] _GEN_1315 = is_Sv39 | state != 2'h0 ? _GEN_1205 : {{24'd0}, pte_addr_r}; // @[tlb.scala 135:37 tlb.scala 47:30]
  ysyx_210539_MaxPeriodFibonacciLFSR_2 select_prng ( // @[PRNG.scala 82:22]
    .clock(select_prng_clock),
    .reset(select_prng_reset),
    .io_out_0(select_prng_io_out_0),
    .io_out_1(select_prng_io_out_1),
    .io_out_2(select_prng_io_out_2),
    .io_out_3(select_prng_io_out_3)
  );
  assign io_va2pa_ready = io_va2pa_vvalid & _T_50 & ~io_flush & ~flush_r; // @[tlb.scala 98:74]
  assign io_va2pa_paddr = out_paddr_r; // @[tlb.scala 113:20]
  assign io_va2pa_pvalid = out_valid_r; // @[tlb.scala 114:21]
  assign io_va2pa_tlb_excep_cause = out_excep_r_cause; // @[tlb.scala 115:24]
  assign io_va2pa_tlb_excep_tval = out_excep_r_tval; // @[tlb.scala 115:24]
  assign io_va2pa_tlb_excep_en = out_excep_r_en; // @[tlb.scala 115:24]
  assign io_dcacheRW_addr = pte_addr_r; // @[tlb.scala 117:22]
  assign io_dcacheRW_wdata = wpte_data_r; // @[tlb.scala 118:23]
  assign io_dcacheRW_dc_mode = dc_mode_r; // @[tlb.scala 119:25]
  assign select_prng_clock = clock;
  assign select_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[tlb.scala 39:26]
      tag_0 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_0 <= _GEN_998;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_1 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_1 <= _GEN_999;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_2 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_2 <= _GEN_1000;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_3 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_3 <= _GEN_1001;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_4 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_4 <= _GEN_1002;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_5 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_5 <= _GEN_1003;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_6 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_6 <= _GEN_1004;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_7 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_7 <= _GEN_1005;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_8 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_8 <= _GEN_1006;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_9 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_9 <= _GEN_1007;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_10 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_10 <= _GEN_1008;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_11 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_11 <= _GEN_1009;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_12 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_12 <= _GEN_1010;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_13 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_13 <= _GEN_1011;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_14 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_14 <= _GEN_1012;
        end
      end
    end
    if (reset) begin // @[tlb.scala 39:26]
      tag_15 <= 52'h0; // @[tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          tag_15 <= _GEN_1013;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_0 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_0 <= _GEN_1030;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_1 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_1 <= _GEN_1031;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_2 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_2 <= _GEN_1032;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_3 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_3 <= _GEN_1033;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_4 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_4 <= _GEN_1034;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_5 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_5 <= _GEN_1035;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_6 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_6 <= _GEN_1036;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_7 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_7 <= _GEN_1037;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_8 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_8 <= _GEN_1038;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_9 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_9 <= _GEN_1039;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_10 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_10 <= _GEN_1040;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_11 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_11 <= _GEN_1041;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_12 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_12 <= _GEN_1042;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_13 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_13 <= _GEN_1043;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_14 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_14 <= _GEN_1044;
        end
      end
    end
    if (reset) begin // @[tlb.scala 40:26]
      paddr_15 <= 20'h0; // @[tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          paddr_15 <= _GEN_1045;
        end
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_0 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_0 <= _GEN_243;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_0 <= _GEN_1078;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_1 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_1 <= _GEN_244;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_1 <= _GEN_1079;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_2 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_2 <= _GEN_245;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_2 <= _GEN_1080;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_3 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_3 <= _GEN_246;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_3 <= _GEN_1081;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_4 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_4 <= _GEN_247;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_4 <= _GEN_1082;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_5 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_5 <= _GEN_248;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_5 <= _GEN_1083;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_6 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_6 <= _GEN_249;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_6 <= _GEN_1084;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_7 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_7 <= _GEN_250;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_7 <= _GEN_1085;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_8 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_8 <= _GEN_251;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_8 <= _GEN_1086;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_9 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_9 <= _GEN_252;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_9 <= _GEN_1087;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_10 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_10 <= _GEN_253;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_10 <= _GEN_1088;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_11 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_11 <= _GEN_254;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_11 <= _GEN_1089;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_12 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_12 <= _GEN_255;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_12 <= _GEN_1090;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_13 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_13 <= _GEN_256;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_13 <= _GEN_1091;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_14 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_14 <= _GEN_257;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_14 <= _GEN_1092;
      end
    end
    if (reset) begin // @[tlb.scala 41:26]
      info_15 <= 10'h0; // @[tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          info_15 <= _GEN_258;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        info_15 <= _GEN_1093;
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_0 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_0 <= _GEN_1046;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_1 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_1 <= _GEN_1047;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_2 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_2 <= _GEN_1048;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_3 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_3 <= _GEN_1049;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_4 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_4 <= _GEN_1050;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_5 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_5 <= _GEN_1051;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_6 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_6 <= _GEN_1052;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_7 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_7 <= _GEN_1053;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_8 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_8 <= _GEN_1054;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_9 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_9 <= _GEN_1055;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_10 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_10 <= _GEN_1056;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_11 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_11 <= _GEN_1057;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_12 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_12 <= _GEN_1058;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_13 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_13 <= _GEN_1059;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_14 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_14 <= _GEN_1060;
        end
      end
    end
    if (reset) begin // @[tlb.scala 42:30]
      pte_addr_15 <= 32'h0; // @[tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_addr_15 <= _GEN_1061;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_0 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_0 <= _GEN_1062;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_1 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_1 <= _GEN_1063;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_2 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_2 <= _GEN_1064;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_3 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_3 <= _GEN_1065;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_4 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_4 <= _GEN_1066;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_5 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_5 <= _GEN_1067;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_6 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_6 <= _GEN_1068;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_7 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_7 <= _GEN_1069;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_8 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_8 <= _GEN_1070;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_9 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_9 <= _GEN_1071;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_10 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_10 <= _GEN_1072;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_11 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_11 <= _GEN_1073;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_12 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_12 <= _GEN_1074;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_13 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_13 <= _GEN_1075;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_14 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_14 <= _GEN_1076;
        end
      end
    end
    if (reset) begin // @[tlb.scala 43:30]
      pte_level_15 <= 2'h0; // @[tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (!(_T_54)) begin // @[Conditional.scala 40:58]
        if (!(_T_68)) begin // @[Conditional.scala 39:67]
          pte_level_15 <= _GEN_1077;
        end
      end
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_0 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_0 <= _GEN_130;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_0 <= _GEN_130;
      end else begin
        valid_0 <= _GEN_1014;
      end
    end else begin
      valid_0 <= _GEN_130;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_1 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_1 <= _GEN_131;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_1 <= _GEN_131;
      end else begin
        valid_1 <= _GEN_1015;
      end
    end else begin
      valid_1 <= _GEN_131;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_2 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_2 <= _GEN_132;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_2 <= _GEN_132;
      end else begin
        valid_2 <= _GEN_1016;
      end
    end else begin
      valid_2 <= _GEN_132;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_3 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_3 <= _GEN_133;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_3 <= _GEN_133;
      end else begin
        valid_3 <= _GEN_1017;
      end
    end else begin
      valid_3 <= _GEN_133;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_4 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_4 <= _GEN_134;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_4 <= _GEN_134;
      end else begin
        valid_4 <= _GEN_1018;
      end
    end else begin
      valid_4 <= _GEN_134;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_5 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_5 <= _GEN_135;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_5 <= _GEN_135;
      end else begin
        valid_5 <= _GEN_1019;
      end
    end else begin
      valid_5 <= _GEN_135;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_6 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_6 <= _GEN_136;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_6 <= _GEN_136;
      end else begin
        valid_6 <= _GEN_1020;
      end
    end else begin
      valid_6 <= _GEN_136;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_7 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_7 <= _GEN_137;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_7 <= _GEN_137;
      end else begin
        valid_7 <= _GEN_1021;
      end
    end else begin
      valid_7 <= _GEN_137;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_8 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_8 <= _GEN_138;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_8 <= _GEN_138;
      end else begin
        valid_8 <= _GEN_1022;
      end
    end else begin
      valid_8 <= _GEN_138;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_9 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_9 <= _GEN_139;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_9 <= _GEN_139;
      end else begin
        valid_9 <= _GEN_1023;
      end
    end else begin
      valid_9 <= _GEN_139;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_10 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_10 <= _GEN_140;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_10 <= _GEN_140;
      end else begin
        valid_10 <= _GEN_1024;
      end
    end else begin
      valid_10 <= _GEN_140;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_11 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_11 <= _GEN_141;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_11 <= _GEN_141;
      end else begin
        valid_11 <= _GEN_1025;
      end
    end else begin
      valid_11 <= _GEN_141;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_12 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_12 <= _GEN_142;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_12 <= _GEN_142;
      end else begin
        valid_12 <= _GEN_1026;
      end
    end else begin
      valid_12 <= _GEN_142;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_13 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_13 <= _GEN_143;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_13 <= _GEN_143;
      end else begin
        valid_13 <= _GEN_1027;
      end
    end else begin
      valid_13 <= _GEN_143;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_14 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_14 <= _GEN_144;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_14 <= _GEN_144;
      end else begin
        valid_14 <= _GEN_1028;
      end
    end else begin
      valid_14 <= _GEN_144;
    end
    if (reset) begin // @[tlb.scala 44:26]
      valid_15 <= 1'h0; // @[tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        valid_15 <= _GEN_145;
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        valid_15 <= _GEN_145;
      end else begin
        valid_15 <= _GEN_1029;
      end
    end else begin
      valid_15 <= _GEN_145;
    end
    if (reset) begin // @[tlb.scala 46:30]
      pre_addr <= 64'h0; // @[tlb.scala 46:30]
    end else if (handshake) begin // @[tlb.scala 101:20]
      pre_addr <= io_va2pa_vaddr; // @[tlb.scala 103:18]
    end else if (io_va2pa_ready & io_va2pa_vvalid) begin // @[tlb.scala 54:44]
      pre_addr <= io_va2pa_vaddr; // @[tlb.scala 55:18]
    end
    if (reset) begin // @[tlb.scala 47:30]
      pte_addr_r <= 32'h0; // @[tlb.scala 47:30]
    end else begin
      pte_addr_r <= _GEN_1315[31:0];
    end
    if (reset) begin // @[tlb.scala 48:30]
      wpte_data_r <= 64'h0; // @[tlb.scala 48:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          wpte_data_r <= _GEN_242;
        end
      end
    end
    if (reset) begin // @[tlb.scala 49:30]
      dc_mode_r <= 5'h0; // @[tlb.scala 49:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (~handshake) begin // @[tlb.scala 139:33]
          dc_mode_r <= 5'h0; // @[tlb.scala 138:27]
        end else begin
          dc_mode_r <= _GEN_261;
        end
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        dc_mode_r <= _GEN_294;
      end else begin
        dc_mode_r <= _GEN_992;
      end
    end
    if (reset) begin // @[tlb.scala 51:30]
      out_valid_r <= 1'h0; // @[tlb.scala 51:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (~handshake) begin // @[tlb.scala 139:33]
          out_valid_r <= _GEN_150;
        end else begin
          out_valid_r <= _GEN_237;
        end
      end else begin
        out_valid_r <= _GEN_150;
      end
    end else begin
      out_valid_r <= io_va2pa_vvalid; // @[tlb.scala 232:21]
    end
    if (reset) begin // @[tlb.scala 52:30]
      out_paddr_r <= 32'h0; // @[tlb.scala 52:30]
    end else begin
      out_paddr_r <= _GEN_1312[31:0];
    end
    if (reset) begin // @[tlb.scala 53:30]
      out_excep_r_cause <= 64'h0; // @[tlb.scala 53:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          out_excep_r_cause <= _GEN_235;
        end
      end
    end
    if (reset) begin // @[tlb.scala 53:30]
      out_excep_r_tval <= 64'h0; // @[tlb.scala 53:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          out_excep_r_tval <= _GEN_236;
        end
      end
    end
    if (reset) begin // @[tlb.scala 53:30]
      out_excep_r_en <= 1'h0; // @[tlb.scala 53:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (~handshake) begin // @[tlb.scala 139:33]
          out_excep_r_en <= _GEN_151;
        end else begin
          out_excep_r_en <= _GEN_234;
        end
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        out_excep_r_en <= _GEN_151;
      end else begin
        out_excep_r_en <= _GEN_996;
      end
    end else begin
      out_excep_r_en <= _GEN_151;
    end
    if (reset) begin // @[tlb.scala 84:24]
      state <= 2'h0; // @[tlb.scala 84:24]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          state <= _GEN_239;
        end
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        state <= _GEN_296;
      end else begin
        state <= _GEN_995;
      end
    end
    if (reset) begin // @[tlb.scala 85:26]
      flush_r <= 1'h0; // @[tlb.scala 85:26]
    end else if (io_flush | flush_r) begin // @[tlb.scala 86:30]
      if (state == 2'h0) begin // @[tlb.scala 87:30]
        flush_r <= 1'h0; // @[tlb.scala 89:21]
      end else begin
        flush_r <= 1'h1; // @[tlb.scala 91:21]
      end
    end
    if (reset) begin // @[tlb.scala 95:27]
      m_type_r <= 2'h0; // @[tlb.scala 95:27]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          m_type_r <= _GEN_260;
        end
      end
    end
    if (reset) begin // @[tlb.scala 130:27]
      select_r <= 4'h0; // @[tlb.scala 130:27]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          select_r <= _GEN_259;
        end
      end
    end
    if (reset) begin // @[tlb.scala 131:26]
      offset <= 8'h0; // @[tlb.scala 131:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          offset <= _GEN_262;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        offset <= _GEN_993;
      end
    end
    if (reset) begin // @[tlb.scala 132:26]
      level <= 2'h0; // @[tlb.scala 132:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          level <= _GEN_263;
        end
      end else if (!(_T_68)) begin // @[Conditional.scala 39:67]
        level <= _GEN_994;
      end
    end
    if (reset) begin // @[tlb.scala 134:28]
      wpte_hs_r <= 1'h0; // @[tlb.scala 134:28]
    end else if (is_Sv39 | state != 2'h0) begin // @[tlb.scala 135:37]
      if (_T_54) begin // @[Conditional.scala 40:58]
        if (!(~handshake)) begin // @[tlb.scala 139:33]
          wpte_hs_r <= _GEN_240;
        end
      end else if (_T_68) begin // @[Conditional.scala 39:67]
        wpte_hs_r <= _GEN_295;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  tag_0 = _RAND_0[51:0];
  _RAND_1 = {2{`RANDOM}};
  tag_1 = _RAND_1[51:0];
  _RAND_2 = {2{`RANDOM}};
  tag_2 = _RAND_2[51:0];
  _RAND_3 = {2{`RANDOM}};
  tag_3 = _RAND_3[51:0];
  _RAND_4 = {2{`RANDOM}};
  tag_4 = _RAND_4[51:0];
  _RAND_5 = {2{`RANDOM}};
  tag_5 = _RAND_5[51:0];
  _RAND_6 = {2{`RANDOM}};
  tag_6 = _RAND_6[51:0];
  _RAND_7 = {2{`RANDOM}};
  tag_7 = _RAND_7[51:0];
  _RAND_8 = {2{`RANDOM}};
  tag_8 = _RAND_8[51:0];
  _RAND_9 = {2{`RANDOM}};
  tag_9 = _RAND_9[51:0];
  _RAND_10 = {2{`RANDOM}};
  tag_10 = _RAND_10[51:0];
  _RAND_11 = {2{`RANDOM}};
  tag_11 = _RAND_11[51:0];
  _RAND_12 = {2{`RANDOM}};
  tag_12 = _RAND_12[51:0];
  _RAND_13 = {2{`RANDOM}};
  tag_13 = _RAND_13[51:0];
  _RAND_14 = {2{`RANDOM}};
  tag_14 = _RAND_14[51:0];
  _RAND_15 = {2{`RANDOM}};
  tag_15 = _RAND_15[51:0];
  _RAND_16 = {1{`RANDOM}};
  paddr_0 = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  paddr_1 = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  paddr_2 = _RAND_18[19:0];
  _RAND_19 = {1{`RANDOM}};
  paddr_3 = _RAND_19[19:0];
  _RAND_20 = {1{`RANDOM}};
  paddr_4 = _RAND_20[19:0];
  _RAND_21 = {1{`RANDOM}};
  paddr_5 = _RAND_21[19:0];
  _RAND_22 = {1{`RANDOM}};
  paddr_6 = _RAND_22[19:0];
  _RAND_23 = {1{`RANDOM}};
  paddr_7 = _RAND_23[19:0];
  _RAND_24 = {1{`RANDOM}};
  paddr_8 = _RAND_24[19:0];
  _RAND_25 = {1{`RANDOM}};
  paddr_9 = _RAND_25[19:0];
  _RAND_26 = {1{`RANDOM}};
  paddr_10 = _RAND_26[19:0];
  _RAND_27 = {1{`RANDOM}};
  paddr_11 = _RAND_27[19:0];
  _RAND_28 = {1{`RANDOM}};
  paddr_12 = _RAND_28[19:0];
  _RAND_29 = {1{`RANDOM}};
  paddr_13 = _RAND_29[19:0];
  _RAND_30 = {1{`RANDOM}};
  paddr_14 = _RAND_30[19:0];
  _RAND_31 = {1{`RANDOM}};
  paddr_15 = _RAND_31[19:0];
  _RAND_32 = {1{`RANDOM}};
  info_0 = _RAND_32[9:0];
  _RAND_33 = {1{`RANDOM}};
  info_1 = _RAND_33[9:0];
  _RAND_34 = {1{`RANDOM}};
  info_2 = _RAND_34[9:0];
  _RAND_35 = {1{`RANDOM}};
  info_3 = _RAND_35[9:0];
  _RAND_36 = {1{`RANDOM}};
  info_4 = _RAND_36[9:0];
  _RAND_37 = {1{`RANDOM}};
  info_5 = _RAND_37[9:0];
  _RAND_38 = {1{`RANDOM}};
  info_6 = _RAND_38[9:0];
  _RAND_39 = {1{`RANDOM}};
  info_7 = _RAND_39[9:0];
  _RAND_40 = {1{`RANDOM}};
  info_8 = _RAND_40[9:0];
  _RAND_41 = {1{`RANDOM}};
  info_9 = _RAND_41[9:0];
  _RAND_42 = {1{`RANDOM}};
  info_10 = _RAND_42[9:0];
  _RAND_43 = {1{`RANDOM}};
  info_11 = _RAND_43[9:0];
  _RAND_44 = {1{`RANDOM}};
  info_12 = _RAND_44[9:0];
  _RAND_45 = {1{`RANDOM}};
  info_13 = _RAND_45[9:0];
  _RAND_46 = {1{`RANDOM}};
  info_14 = _RAND_46[9:0];
  _RAND_47 = {1{`RANDOM}};
  info_15 = _RAND_47[9:0];
  _RAND_48 = {1{`RANDOM}};
  pte_addr_0 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  pte_addr_1 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  pte_addr_2 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  pte_addr_3 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  pte_addr_4 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  pte_addr_5 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  pte_addr_6 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  pte_addr_7 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  pte_addr_8 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  pte_addr_9 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  pte_addr_10 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  pte_addr_11 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  pte_addr_12 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  pte_addr_13 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  pte_addr_14 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  pte_addr_15 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  pte_level_0 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  pte_level_1 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  pte_level_2 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  pte_level_3 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  pte_level_4 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  pte_level_5 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  pte_level_6 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  pte_level_7 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  pte_level_8 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  pte_level_9 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  pte_level_10 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  pte_level_11 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  pte_level_12 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  pte_level_13 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  pte_level_14 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  pte_level_15 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  valid_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_4 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_5 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_6 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_7 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_8 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_9 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_10 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_11 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_12 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_13 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_14 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_15 = _RAND_95[0:0];
  _RAND_96 = {2{`RANDOM}};
  pre_addr = _RAND_96[63:0];
  _RAND_97 = {1{`RANDOM}};
  pte_addr_r = _RAND_97[31:0];
  _RAND_98 = {2{`RANDOM}};
  wpte_data_r = _RAND_98[63:0];
  _RAND_99 = {1{`RANDOM}};
  dc_mode_r = _RAND_99[4:0];
  _RAND_100 = {1{`RANDOM}};
  out_valid_r = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  out_paddr_r = _RAND_101[31:0];
  _RAND_102 = {2{`RANDOM}};
  out_excep_r_cause = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  out_excep_r_tval = _RAND_103[63:0];
  _RAND_104 = {1{`RANDOM}};
  out_excep_r_en = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  state = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  flush_r = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  m_type_r = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  select_r = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  offset = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  level = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  wpte_hs_r = _RAND_111[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_DcacheSelector(
  input         clock,
  input         reset,
  input  [31:0] io_tlb_if2dc_addr,
  output [63:0] io_tlb_if2dc_rdata,
  output        io_tlb_if2dc_rvalid,
  input  [63:0] io_tlb_if2dc_wdata,
  input  [4:0]  io_tlb_if2dc_dc_mode,
  output        io_tlb_if2dc_ready,
  input  [31:0] io_tlb_mem2dc_addr,
  output [63:0] io_tlb_mem2dc_rdata,
  output        io_tlb_mem2dc_rvalid,
  input  [63:0] io_tlb_mem2dc_wdata,
  input  [4:0]  io_tlb_mem2dc_dc_mode,
  output        io_tlb_mem2dc_ready,
  input  [31:0] io_mem2dc_addr,
  output [63:0] io_mem2dc_rdata,
  output        io_mem2dc_rvalid,
  input  [63:0] io_mem2dc_wdata,
  input  [4:0]  io_mem2dc_dc_mode,
  input  [4:0]  io_mem2dc_amo,
  output        io_mem2dc_ready,
  input  [31:0] io_dma2dc_addr,
  output [63:0] io_dma2dc_rdata,
  output        io_dma2dc_rvalid,
  input  [63:0] io_dma2dc_wdata,
  input  [4:0]  io_dma2dc_dc_mode,
  output        io_dma2dc_ready,
  output [31:0] io_select_addr,
  input  [63:0] io_select_rdata,
  input         io_select_rvalid,
  output [63:0] io_select_wdata,
  output [4:0]  io_select_dc_mode,
  output [4:0]  io_select_amo,
  input         io_select_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] pre_idx; // @[dcache.scala 30:26]
  reg  busy; // @[dcache.scala 31:26]
  wire  _GEN_0 = io_select_rvalid ? 1'h0 : busy; // @[dcache.scala 37:27 dcache.scala 38:14 dcache.scala 31:26]
  wire [1:0] _GEN_1 = io_dma2dc_dc_mode != 5'h0 ? 2'h3 : pre_idx; // @[dcache.scala 65:47 dcache.scala 66:17 dcache.scala 30:26]
  wire  _GEN_2 = io_dma2dc_dc_mode != 5'h0 ? io_select_ready : _GEN_0; // @[dcache.scala 65:47 dcache.scala 67:17]
  wire [31:0] _GEN_3 = io_dma2dc_dc_mode != 5'h0 ? io_dma2dc_addr : 32'h0; // @[dcache.scala 65:47 dcache.scala 68:29 dcache.scala 32:25]
  wire [63:0] _GEN_4 = io_dma2dc_dc_mode != 5'h0 ? io_dma2dc_wdata : 64'h0; // @[dcache.scala 65:47 dcache.scala 69:29 dcache.scala 33:25]
  wire [4:0] _GEN_5 = io_dma2dc_dc_mode != 5'h0 ? io_dma2dc_dc_mode : 5'h0; // @[dcache.scala 65:47 dcache.scala 70:29 dcache.scala 34:25]
  wire  _GEN_7 = io_dma2dc_dc_mode != 5'h0 & io_select_ready; // @[dcache.scala 65:47 dcache.scala 72:29 dcache.scala 29:69]
  wire [1:0] _GEN_8 = io_tlb_if2dc_dc_mode != 5'h0 ? 2'h2 : _GEN_1; // @[dcache.scala 57:50 dcache.scala 58:17]
  wire  _GEN_9 = io_tlb_if2dc_dc_mode != 5'h0 ? io_select_ready : _GEN_2; // @[dcache.scala 57:50 dcache.scala 59:17]
  wire [31:0] _GEN_10 = io_tlb_if2dc_dc_mode != 5'h0 ? io_tlb_if2dc_addr : _GEN_3; // @[dcache.scala 57:50 dcache.scala 60:29]
  wire [63:0] _GEN_11 = io_tlb_if2dc_dc_mode != 5'h0 ? io_tlb_if2dc_wdata : _GEN_4; // @[dcache.scala 57:50 dcache.scala 61:29]
  wire [4:0] _GEN_12 = io_tlb_if2dc_dc_mode != 5'h0 ? io_tlb_if2dc_dc_mode : _GEN_5; // @[dcache.scala 57:50 dcache.scala 62:29]
  wire  _GEN_14 = io_tlb_if2dc_dc_mode != 5'h0 & io_select_ready; // @[dcache.scala 57:50 dcache.scala 64:29 dcache.scala 23:69]
  wire  _GEN_15 = io_tlb_if2dc_dc_mode != 5'h0 ? 1'h0 : _GEN_7; // @[dcache.scala 57:50 dcache.scala 29:69]
  wire [31:0] _GEN_18 = io_tlb_mem2dc_dc_mode != 5'h0 ? io_tlb_mem2dc_addr : _GEN_10; // @[dcache.scala 49:51 dcache.scala 52:29]
  wire [63:0] _GEN_19 = io_tlb_mem2dc_dc_mode != 5'h0 ? io_tlb_mem2dc_wdata : _GEN_11; // @[dcache.scala 49:51 dcache.scala 53:29]
  wire [4:0] _GEN_20 = io_tlb_mem2dc_dc_mode != 5'h0 ? io_tlb_mem2dc_dc_mode : _GEN_12; // @[dcache.scala 49:51 dcache.scala 54:29]
  wire  _GEN_22 = io_tlb_mem2dc_dc_mode != 5'h0 & io_select_ready; // @[dcache.scala 49:51 dcache.scala 56:29 dcache.scala 25:69]
  wire  _GEN_23 = io_tlb_mem2dc_dc_mode != 5'h0 ? 1'h0 : _GEN_14; // @[dcache.scala 49:51 dcache.scala 23:69]
  wire  _GEN_24 = io_tlb_mem2dc_dc_mode != 5'h0 ? 1'h0 : _GEN_15; // @[dcache.scala 49:51 dcache.scala 29:69]
  wire [31:0] _GEN_27 = io_mem2dc_dc_mode != 5'h0 ? io_mem2dc_addr : _GEN_18; // @[dcache.scala 41:47 dcache.scala 44:29]
  wire [63:0] _GEN_28 = io_mem2dc_dc_mode != 5'h0 ? io_mem2dc_wdata : _GEN_19; // @[dcache.scala 41:47 dcache.scala 45:29]
  wire [4:0] _GEN_29 = io_mem2dc_dc_mode != 5'h0 ? io_mem2dc_dc_mode : _GEN_20; // @[dcache.scala 41:47 dcache.scala 46:29]
  wire [4:0] _GEN_30 = io_mem2dc_dc_mode != 5'h0 ? io_mem2dc_amo : 5'h0; // @[dcache.scala 41:47 dcache.scala 47:29]
  wire  _GEN_31 = io_mem2dc_dc_mode != 5'h0 & io_select_ready; // @[dcache.scala 41:47 dcache.scala 48:29 dcache.scala 36:25]
  wire  _GEN_32 = io_mem2dc_dc_mode != 5'h0 ? 1'h0 : _GEN_22; // @[dcache.scala 41:47 dcache.scala 25:69]
  wire  _GEN_33 = io_mem2dc_dc_mode != 5'h0 ? 1'h0 : _GEN_23; // @[dcache.scala 41:47 dcache.scala 23:69]
  wire  _GEN_34 = io_mem2dc_dc_mode != 5'h0 ? 1'h0 : _GEN_24; // @[dcache.scala 41:47 dcache.scala 29:69]
  assign io_tlb_if2dc_rdata = io_select_rdata; // @[dcache.scala 22:29]
  assign io_tlb_if2dc_rvalid = io_select_rvalid & pre_idx == 2'h2; // @[dcache.scala 76:49]
  assign io_tlb_if2dc_ready = busy & ~io_select_rvalid ? 1'h0 : _GEN_33; // @[dcache.scala 40:36 dcache.scala 23:69]
  assign io_tlb_mem2dc_rdata = io_select_rdata; // @[dcache.scala 24:29]
  assign io_tlb_mem2dc_rvalid = io_select_rvalid & pre_idx == 2'h1; // @[dcache.scala 75:49]
  assign io_tlb_mem2dc_ready = busy & ~io_select_rvalid ? 1'h0 : _GEN_32; // @[dcache.scala 40:36 dcache.scala 25:69]
  assign io_mem2dc_rdata = io_select_rdata; // @[dcache.scala 26:29]
  assign io_mem2dc_rvalid = io_select_rvalid & pre_idx == 2'h0; // @[dcache.scala 74:49]
  assign io_mem2dc_ready = busy & ~io_select_rvalid ? 1'h0 : _GEN_31; // @[dcache.scala 40:36 dcache.scala 36:25]
  assign io_dma2dc_rdata = io_select_rdata; // @[dcache.scala 28:29]
  assign io_dma2dc_rvalid = io_select_rvalid & pre_idx == 2'h3; // @[dcache.scala 77:49]
  assign io_dma2dc_ready = busy & ~io_select_rvalid ? 1'h0 : _GEN_34; // @[dcache.scala 40:36 dcache.scala 29:69]
  assign io_select_addr = busy & ~io_select_rvalid ? 32'h0 : _GEN_27; // @[dcache.scala 40:36 dcache.scala 32:25]
  assign io_select_wdata = busy & ~io_select_rvalid ? 64'h0 : _GEN_28; // @[dcache.scala 40:36 dcache.scala 33:25]
  assign io_select_dc_mode = busy & ~io_select_rvalid ? 5'h0 : _GEN_29; // @[dcache.scala 40:36 dcache.scala 34:25]
  assign io_select_amo = busy & ~io_select_rvalid ? 5'h0 : _GEN_30; // @[dcache.scala 40:36 dcache.scala 35:25]
  always @(posedge clock) begin
    if (reset) begin // @[dcache.scala 30:26]
      pre_idx <= 2'h0; // @[dcache.scala 30:26]
    end else if (!(busy & ~io_select_rvalid)) begin // @[dcache.scala 40:36]
      if (io_mem2dc_dc_mode != 5'h0) begin // @[dcache.scala 41:47]
        pre_idx <= 2'h0; // @[dcache.scala 42:17]
      end else if (io_tlb_mem2dc_dc_mode != 5'h0) begin // @[dcache.scala 49:51]
        pre_idx <= 2'h1; // @[dcache.scala 50:17]
      end else begin
        pre_idx <= _GEN_8;
      end
    end
    if (reset) begin // @[dcache.scala 31:26]
      busy <= 1'h0; // @[dcache.scala 31:26]
    end else if (busy & ~io_select_rvalid) begin // @[dcache.scala 40:36]
      if (io_select_rvalid) begin // @[dcache.scala 37:27]
        busy <= 1'h0; // @[dcache.scala 38:14]
      end
    end else if (io_mem2dc_dc_mode != 5'h0) begin // @[dcache.scala 41:47]
      busy <= io_select_ready; // @[dcache.scala 43:17]
    end else if (io_tlb_mem2dc_dc_mode != 5'h0) begin // @[dcache.scala 49:51]
      busy <= io_select_ready; // @[dcache.scala 51:17]
    end else begin
      busy <= _GEN_9;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pre_idx = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  busy = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_CLINT(
  input         clock,
  input         reset,
  input  [31:0] io_rw_addr,
  output [63:0] io_rw_rdata,
  input  [63:0] io_rw_wdata,
  input         io_rw_wvalid,
  output        io_intr_raise,
  output        io_intr_clear,
  output        io_intr_msip_raise,
  output        io_intr_msip_clear
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtime; // @[clint.scala 21:24]
  reg [63:0] mtimecmp; // @[clint.scala 22:27]
  reg [63:0] ipi; // @[clint.scala 23:22]
  reg [1:0] count; // @[clint.scala 24:24]
  reg  clear_r; // @[clint.scala 25:26]
  wire [1:0] _count_T_1 = count + 2'h1; // @[clint.scala 27:20]
  wire [63:0] _mtime_T_1 = mtime + 64'h1; // @[clint.scala 29:24]
  wire [63:0] _GEN_0 = count == 2'h0 ? _mtime_T_1 : mtime; // @[clint.scala 28:24 clint.scala 29:15 clint.scala 21:24]
  wire [63:0] _GEN_2 = io_rw_addr == 32'h200bff8 ? mtime : 64'h0; // @[clint.scala 35:31 clint.scala 36:24 clint.scala 34:17]
  wire [63:0] _GEN_6 = io_rw_addr == 32'h2004000 ? mtimecmp : _GEN_2; // @[clint.scala 41:34 clint.scala 42:24]
  wire  _GEN_8 = io_rw_addr == 32'h2004000 & io_rw_wvalid; // @[clint.scala 41:34 clint.scala 26:13]
  wire  _GEN_10 = io_rw_wvalid & io_rw_wdata[0]; // @[clint.scala 50:27 clint.scala 52:32 clint.scala 33:20]
  wire  _GEN_11 = io_rw_wvalid & ~io_rw_wdata[0]; // @[clint.scala 50:27 clint.scala 53:32 clint.scala 33:20]
  assign io_rw_rdata = io_rw_addr == 32'h2000000 ? ipi : _GEN_6; // @[clint.scala 48:29 clint.scala 49:24]
  assign io_intr_raise = mtime > mtimecmp; // @[clint.scala 31:28]
  assign io_intr_clear = clear_r; // @[clint.scala 32:19]
  assign io_intr_msip_raise = io_rw_addr == 32'h2000000 & _GEN_10; // @[clint.scala 48:29 clint.scala 33:20]
  assign io_intr_msip_clear = io_rw_addr == 32'h2000000 & _GEN_11; // @[clint.scala 48:29 clint.scala 33:20]
  always @(posedge clock) begin
    if (reset) begin // @[clint.scala 21:24]
      mtime <= 64'h0; // @[clint.scala 21:24]
    end else if (io_rw_addr == 32'h200bff8) begin // @[clint.scala 35:31]
      if (io_rw_wvalid) begin // @[clint.scala 37:27]
        mtime <= io_rw_wdata; // @[clint.scala 38:19]
      end else begin
        mtime <= _GEN_0;
      end
    end else begin
      mtime <= _GEN_0;
    end
    if (reset) begin // @[clint.scala 22:27]
      mtimecmp <= 64'h0; // @[clint.scala 22:27]
    end else if (io_rw_addr == 32'h2004000) begin // @[clint.scala 41:34]
      if (io_rw_wvalid) begin // @[clint.scala 43:27]
        mtimecmp <= io_rw_wdata; // @[clint.scala 44:22]
      end
    end
    if (reset) begin // @[clint.scala 23:22]
      ipi <= 64'h0; // @[clint.scala 23:22]
    end else if (io_rw_addr == 32'h2000000) begin // @[clint.scala 48:29]
      if (io_rw_wvalid) begin // @[clint.scala 50:27]
        ipi <= io_rw_wdata; // @[clint.scala 51:17]
      end
    end
    if (reset) begin // @[clint.scala 24:24]
      count <= 2'h0; // @[clint.scala 24:24]
    end else begin
      count <= _count_T_1; // @[clint.scala 27:11]
    end
    if (reset) begin // @[clint.scala 25:26]
      clear_r <= 1'h0; // @[clint.scala 25:26]
    end else begin
      clear_r <= _GEN_8;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtime = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtimecmp = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  ipi = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  count = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  clear_r = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_Plic(
  input         clock,
  input         reset,
  input         io_intr_in1,
  output        io_intr_out_m_raise,
  output        io_intr_out_m_clear,
  output        io_intr_out_s_raise,
  output        io_intr_out_s_clear,
  input  [31:0] io_rw_addr,
  output [63:0] io_rw_rdata,
  input  [63:0] io_rw_wdata,
  input         io_rw_wvalid,
  input         io_rw_arvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] priority_; // @[plic.scala 34:27]
  reg [31:0] pending; // @[plic.scala 35:26]
  reg [31:0] intr_enable1; // @[plic.scala 36:31]
  reg [31:0] intr_enable2; // @[plic.scala 37:31]
  reg [31:0] threshold1; // @[plic.scala 38:29]
  reg [31:0] threshold2; // @[plic.scala 39:29]
  reg [31:0] claim1; // @[plic.scala 40:25]
  reg [31:0] claim2; // @[plic.scala 41:25]
  reg  clear_r; // @[plic.scala 43:26]
  wire [63:0] _GEN_32 = {{32'd0}, pending}; // @[plic.scala 23:18]
  wire [63:0] _pending_T_1 = _GEN_32 & 64'hfffffffffffffffd; // @[plic.scala 23:18]
  wire [63:0] _pending_T_4 = _pending_T_1 | 64'h2; // @[plic.scala 23:27]
  wire [63:0] _GEN_0 = io_intr_in1 ? _pending_T_4 : {{32'd0}, pending}; // @[plic.scala 51:22 plic.scala 52:17 plic.scala 35:26]
  wire [31:0] _GEN_1 = io_intr_out_m_raise ? 32'h1 : claim1; // @[plic.scala 54:30 plic.scala 55:16 plic.scala 40:25]
  wire [31:0] _GEN_2 = io_intr_out_s_raise ? 32'h1 : claim2; // @[plic.scala 57:30 plic.scala 58:16 plic.scala 41:25]
  wire [63:0] _GEN_3 = io_rw_wvalid ? io_rw_wdata : {{32'd0}, priority_}; // @[plic.scala 63:27 plic.scala 64:22 plic.scala 34:27]
  wire [31:0] _GEN_4 = io_rw_addr == 32'hc000004 ? priority_ : 32'h0; // @[plic.scala 61:39 plic.scala 62:21 plic.scala 50:17]
  wire [63:0] _GEN_5 = io_rw_addr == 32'hc000004 ? _GEN_3 : {{32'd0}, priority_}; // @[plic.scala 61:39 plic.scala 34:27]
  wire [63:0] _GEN_6 = io_rw_wvalid ? io_rw_wdata : {{32'd0}, intr_enable1}; // @[plic.scala 69:27 plic.scala 70:26 plic.scala 36:31]
  wire [31:0] _GEN_7 = io_rw_addr == 32'hc002000 ? intr_enable1 : _GEN_4; // @[plic.scala 67:38 plic.scala 68:21]
  wire [63:0] _GEN_8 = io_rw_addr == 32'hc002000 ? _GEN_6 : {{32'd0}, intr_enable1}; // @[plic.scala 67:38 plic.scala 36:31]
  wire [63:0] _GEN_9 = io_rw_wvalid ? io_rw_wdata : {{32'd0}, intr_enable2}; // @[plic.scala 75:27 plic.scala 76:26 plic.scala 37:31]
  wire [31:0] _GEN_10 = io_rw_addr == 32'hc002100 ? intr_enable2 : _GEN_7; // @[plic.scala 73:38 plic.scala 74:21]
  wire [63:0] _GEN_11 = io_rw_addr == 32'hc002100 ? _GEN_9 : {{32'd0}, intr_enable2}; // @[plic.scala 73:38 plic.scala 37:31]
  wire [5:0] pending_bit_idx = claim1[5:0]; // @[plic.scala 21:26]
  wire [63:0] pending_mask_1 = 64'h1 << pending_bit_idx; // @[plic.scala 22:24]
  wire [63:0] _pending_T_5 = ~pending_mask_1; // @[plic.scala 23:20]
  wire [63:0] _pending_T_6 = _GEN_32 & _pending_T_5; // @[plic.scala 23:18]
  wire [63:0] _pending_T_7 = 64'h0 << pending_bit_idx; // @[plic.scala 23:37]
  wire [63:0] _pending_T_8 = _pending_T_7 & pending_mask_1; // @[plic.scala 23:49]
  wire [63:0] _pending_T_9 = _pending_T_6 | _pending_T_8; // @[plic.scala 23:27]
  wire [63:0] _GEN_12 = io_rw_arvalid ? _pending_T_9 : _GEN_0; // @[plic.scala 81:28 plic.scala 82:21]
  wire [31:0] _GEN_15 = io_rw_addr == 32'hc200004 ? claim1 : _GEN_10; // @[plic.scala 79:37 plic.scala 80:21]
  wire [63:0] _GEN_16 = io_rw_addr == 32'hc200004 ? _GEN_12 : _GEN_0; // @[plic.scala 79:37]
  wire  _GEN_17 = io_rw_addr == 32'hc200004 & io_rw_arvalid; // @[plic.scala 79:37 plic.scala 44:13]
  wire [5:0] pending_bit_idx_1 = claim2[5:0]; // @[plic.scala 21:26]
  wire [63:0] pending_mask_2 = 64'h1 << pending_bit_idx_1; // @[plic.scala 22:24]
  wire [63:0] _pending_T_10 = ~pending_mask_2; // @[plic.scala 23:20]
  wire [63:0] _pending_T_11 = _GEN_32 & _pending_T_10; // @[plic.scala 23:18]
  wire [63:0] _pending_T_12 = 64'h0 << pending_bit_idx_1; // @[plic.scala 23:37]
  wire [63:0] _pending_T_13 = _pending_T_12 & pending_mask_2; // @[plic.scala 23:49]
  wire [63:0] _pending_T_14 = _pending_T_11 | _pending_T_13; // @[plic.scala 23:27]
  wire [63:0] _GEN_19 = io_rw_arvalid ? _pending_T_14 : _GEN_16; // @[plic.scala 91:28 plic.scala 92:21]
  wire  _GEN_20 = io_rw_arvalid | _GEN_17; // @[plic.scala 91:28 plic.scala 93:21]
  wire [31:0] _GEN_22 = io_rw_addr == 32'hc201004 ? claim2 : _GEN_15; // @[plic.scala 89:37 plic.scala 90:21]
  wire [63:0] _GEN_23 = io_rw_addr == 32'hc201004 ? _GEN_19 : _GEN_16; // @[plic.scala 89:37]
  wire [63:0] _GEN_26 = io_rw_wvalid ? io_rw_wdata : {{32'd0}, threshold1}; // @[plic.scala 101:27 plic.scala 102:24 plic.scala 38:29]
  wire [31:0] _GEN_27 = io_rw_addr == 32'hc200000 ? threshold1 : _GEN_22; // @[plic.scala 99:41 plic.scala 100:21]
  wire [63:0] _GEN_28 = io_rw_addr == 32'hc200000 ? _GEN_26 : {{32'd0}, threshold1}; // @[plic.scala 99:41 plic.scala 38:29]
  wire [63:0] _GEN_29 = io_rw_wvalid ? io_rw_wdata : {{32'd0}, threshold2}; // @[plic.scala 107:27 plic.scala 108:24 plic.scala 39:29]
  wire [31:0] _GEN_30 = io_rw_addr == 32'hc201000 ? threshold2 : _GEN_27; // @[plic.scala 105:41 plic.scala 106:21]
  wire [63:0] _GEN_31 = io_rw_addr == 32'hc201000 ? _GEN_29 : {{32'd0}, threshold2}; // @[plic.scala 105:41 plic.scala 39:29]
  assign io_intr_out_m_raise = pending[1] & priority_ >= threshold1; // @[plic.scala 48:39]
  assign io_intr_out_m_clear = clear_r; // @[plic.scala 49:25]
  assign io_intr_out_s_raise = pending[1] & priority_ >= threshold2; // @[plic.scala 46:39]
  assign io_intr_out_s_clear = clear_r; // @[plic.scala 47:25]
  assign io_rw_rdata = {{32'd0}, _GEN_30}; // @[plic.scala 105:41 plic.scala 106:21]
  always @(posedge clock) begin
    if (reset) begin // @[plic.scala 34:27]
      priority_ <= 32'h0; // @[plic.scala 34:27]
    end else begin
      priority_ <= _GEN_5[31:0];
    end
    if (reset) begin // @[plic.scala 35:26]
      pending <= 32'h0; // @[plic.scala 35:26]
    end else begin
      pending <= _GEN_23[31:0];
    end
    if (reset) begin // @[plic.scala 36:31]
      intr_enable1 <= 32'h0; // @[plic.scala 36:31]
    end else begin
      intr_enable1 <= _GEN_8[31:0];
    end
    if (reset) begin // @[plic.scala 37:31]
      intr_enable2 <= 32'h0; // @[plic.scala 37:31]
    end else begin
      intr_enable2 <= _GEN_11[31:0];
    end
    if (reset) begin // @[plic.scala 38:29]
      threshold1 <= 32'h0; // @[plic.scala 38:29]
    end else begin
      threshold1 <= _GEN_28[31:0];
    end
    if (reset) begin // @[plic.scala 39:29]
      threshold2 <= 32'h0; // @[plic.scala 39:29]
    end else begin
      threshold2 <= _GEN_31[31:0];
    end
    if (reset) begin // @[plic.scala 40:25]
      claim1 <= 32'h0; // @[plic.scala 40:25]
    end else if (io_rw_addr == 32'hc200004) begin // @[plic.scala 79:37]
      if (io_rw_arvalid) begin // @[plic.scala 81:28]
        claim1 <= 32'h0; // @[plic.scala 84:20]
      end else begin
        claim1 <= _GEN_1;
      end
    end else begin
      claim1 <= _GEN_1;
    end
    if (reset) begin // @[plic.scala 41:25]
      claim2 <= 32'h0; // @[plic.scala 41:25]
    end else if (io_rw_addr == 32'hc201004) begin // @[plic.scala 89:37]
      if (io_rw_arvalid) begin // @[plic.scala 91:28]
        claim2 <= 32'h0; // @[plic.scala 94:20]
      end else begin
        claim2 <= _GEN_2;
      end
    end else begin
      claim2 <= _GEN_2;
    end
    if (reset) begin // @[plic.scala 43:26]
      clear_r <= 1'h0; // @[plic.scala 43:26]
    end else if (io_rw_addr == 32'hc201004) begin // @[plic.scala 89:37]
      clear_r <= _GEN_20;
    end else begin
      clear_r <= _GEN_17;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  priority_ = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  pending = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  intr_enable1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  intr_enable2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  threshold1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  threshold2 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  claim1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  claim2 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  clear_r = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210539_DmaBridge(
  input         clock,
  input         reset,
  output        io_dmaAxi_awready,
  input         io_dmaAxi_awvalid,
  input  [31:0] io_dmaAxi_awaddr,
  input  [3:0]  io_dmaAxi_awid,
  input  [7:0]  io_dmaAxi_awlen,
  input  [2:0]  io_dmaAxi_awsize,
  output        io_dmaAxi_wready,
  input         io_dmaAxi_wvalid,
  input  [63:0] io_dmaAxi_wdata,
  input  [7:0]  io_dmaAxi_wstrb,
  input         io_dmaAxi_bready,
  output        io_dmaAxi_bvalid,
  output [3:0]  io_dmaAxi_bid,
  output        io_dmaAxi_arready,
  input         io_dmaAxi_arvalid,
  input  [31:0] io_dmaAxi_araddr,
  input  [3:0]  io_dmaAxi_arid,
  input  [7:0]  io_dmaAxi_arlen,
  input  [2:0]  io_dmaAxi_arsize,
  input         io_dmaAxi_rready,
  output        io_dmaAxi_rvalid,
  output [63:0] io_dmaAxi_rdata,
  output        io_dmaAxi_rlast,
  output [3:0]  io_dmaAxi_rid,
  output [31:0] io_dcRW_addr,
  input  [63:0] io_dcRW_rdata,
  input         io_dcRW_rvalid,
  output [63:0] io_dcRW_wdata,
  output [4:0]  io_dcRW_dc_mode,
  input         io_dcRW_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[dma.scala 18:24]
  reg  awready_r; // @[dma.scala 20:30]
  reg  wready_r; // @[dma.scala 21:30]
  reg  bvalid_r; // @[dma.scala 22:30]
  reg [3:0] bid_r; // @[dma.scala 24:30]
  reg  arready_r; // @[dma.scala 25:30]
  reg  rvalid_r; // @[dma.scala 26:30]
  reg [63:0] rdata_r; // @[dma.scala 28:30]
  reg  rlast_r; // @[dma.scala 29:30]
  reg [3:0] rid_r; // @[dma.scala 30:30]
  reg [31:0] dc_addr_r; // @[dma.scala 32:30]
  reg [63:0] dc_wdata_r; // @[dma.scala 33:30]
  reg [4:0] dc_mode_r; // @[dma.scala 34:30]
  reg [63:0] data_buf_r; // @[dma.scala 35:30]
  reg [7:0] data_strb_r; // @[dma.scala 36:30]
  reg [31:0] addr_r; // @[dma.scala 39:30]
  reg [3:0] id_r; // @[dma.scala 40:30]
  reg [7:0] len_r; // @[dma.scala 41:30]
  reg [7:0] size_r; // @[dma.scala 42:30]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _GEN_1 = io_dmaAxi_arvalid | arready_r; // @[dma.scala 48:36 dma.scala 50:29 dma.scala 25:30]
  wire  _GEN_3 = io_dmaAxi_awvalid | awready_r; // @[dma.scala 52:36 dma.scala 54:29 dma.scala 20:30]
  wire  _T_1 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire [7:0] _size_r_T = 8'h1 << io_dmaAxi_arsize; // @[dma.scala 62:32]
  wire [31:0] _dc_addr_r_T_1 = io_dmaAxi_araddr & 32'hfffffff8; // @[dma.scala 65:45]
  wire  _T_2 = 3'h6 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = io_dcRW_ready & dc_mode_r != 5'h0; // @[dma.scala 69:32]
  wire [4:0] _GEN_4 = io_dcRW_ready & dc_mode_r != 5'h0 ? 5'h0 : dc_mode_r; // @[dma.scala 69:60 dma.scala 70:27 dma.scala 34:30]
  wire [63:0] _GEN_5 = io_dcRW_rvalid ? io_dcRW_rdata : data_buf_r; // @[dma.scala 72:33 dma.scala 73:28 dma.scala 35:30]
  wire [2:0] _GEN_6 = io_dcRW_rvalid ? 3'h2 : state; // @[dma.scala 72:33 dma.scala 74:23 dma.scala 18:24]
  wire  _T_5 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _rlast_r_T = len_r == 8'h0; // @[dma.scala 80:30]
  wire [7:0] _len_r_T_1 = len_r - 8'h1; // @[dma.scala 88:36]
  wire [31:0] _GEN_190 = {{24'd0}, size_r}; // @[dma.scala 89:42]
  wire [31:0] _dc_addr_r_T_3 = addr_r + _GEN_190; // @[dma.scala 89:42]
  wire [31:0] _dc_addr_r_T_5 = _dc_addr_r_T_3 & 32'hfffffff8; // @[dma.scala 89:52]
  wire [2:0] _GEN_7 = rlast_r ? 3'h0 : 3'h6; // @[dma.scala 85:30 dma.scala 86:27 dma.scala 92:27]
  wire [7:0] _GEN_8 = rlast_r ? len_r : _len_r_T_1; // @[dma.scala 85:30 dma.scala 41:30 dma.scala 88:27]
  wire [31:0] _GEN_9 = rlast_r ? dc_addr_r : _dc_addr_r_T_5; // @[dma.scala 85:30 dma.scala 32:30 dma.scala 89:31]
  wire [31:0] _GEN_10 = rlast_r ? addr_r : _dc_addr_r_T_3; // @[dma.scala 85:30 dma.scala 39:30 dma.scala 90:28]
  wire [4:0] _GEN_11 = rlast_r ? dc_mode_r : 5'h7; // @[dma.scala 85:30 dma.scala 34:30 dma.scala 91:31]
  wire  _GEN_12 = io_dmaAxi_rready & rvalid_r ? 1'h0 : 1'h1; // @[dma.scala 83:47 dma.scala 84:26 dma.scala 79:22]
  wire [2:0] _GEN_13 = io_dmaAxi_rready & rvalid_r ? _GEN_7 : state; // @[dma.scala 83:47 dma.scala 18:24]
  wire [7:0] _GEN_14 = io_dmaAxi_rready & rvalid_r ? _GEN_8 : len_r; // @[dma.scala 83:47 dma.scala 41:30]
  wire [31:0] _GEN_15 = io_dmaAxi_rready & rvalid_r ? _GEN_9 : dc_addr_r; // @[dma.scala 83:47 dma.scala 32:30]
  wire [31:0] _GEN_16 = io_dmaAxi_rready & rvalid_r ? _GEN_10 : addr_r; // @[dma.scala 83:47 dma.scala 39:30]
  wire [4:0] _GEN_17 = io_dmaAxi_rready & rvalid_r ? _GEN_11 : dc_mode_r; // @[dma.scala 83:47 dma.scala 34:30]
  wire  _T_7 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire [31:0] _dc_addr_r_T_7 = io_dmaAxi_awaddr & 32'hfffffff8; // @[dma.scala 99:45]
  wire [7:0] _size_r_T_1 = 8'h1 << io_dmaAxi_awsize; // @[dma.scala 102:32]
  wire  _T_8 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _GEN_18 = io_dmaAxi_wvalid & wready_r ? 1'h0 : wready_r; // @[dma.scala 108:47 dma.scala 109:29 dma.scala 21:30]
  wire [63:0] _GEN_19 = io_dmaAxi_wvalid & wready_r ? io_dmaAxi_wdata : data_buf_r; // @[dma.scala 108:47 dma.scala 110:29 dma.scala 35:30]
  wire [7:0] _GEN_20 = io_dmaAxi_wvalid & wready_r ? io_dmaAxi_wstrb : data_strb_r; // @[dma.scala 108:47 dma.scala 111:29 dma.scala 36:30]
  wire [2:0] _GEN_22 = io_dmaAxi_wvalid & wready_r ? 3'h7 : state; // @[dma.scala 108:47 dma.scala 113:29 dma.scala 18:24]
  wire  _T_10 = 3'h7 == state; // @[Conditional.scala 37:30]
  wire  _GEN_23 = _rlast_r_T | bvalid_r; // @[dma.scala 120:36 dma.scala 121:30 dma.scala 22:30]
  wire [3:0] _GEN_25 = _rlast_r_T ? id_r : bid_r; // @[dma.scala 120:36 dma.scala 123:29 dma.scala 24:30]
  wire [2:0] _GEN_26 = _rlast_r_T ? 3'h5 : 3'h4; // @[dma.scala 120:36 dma.scala 124:29 dma.scala 126:27]
  wire  _GEN_27 = _rlast_r_T ? wready_r : 1'h1; // @[dma.scala 120:36 dma.scala 21:30 dma.scala 127:30]
  wire [7:0] _GEN_28 = _rlast_r_T ? len_r : _len_r_T_1; // @[dma.scala 120:36 dma.scala 41:30 dma.scala 128:27]
  wire [7:0] _data_strb_r_T = {{1'd0}, data_strb_r[7:1]}; // @[dma.scala 135:48]
  wire [63:0] _data_buf_r_T = {{8'd0}, data_buf_r[63:8]}; // @[dma.scala 136:47]
  wire [31:0] _dc_addr_r_T_13 = dc_addr_r + 32'h1; // @[dma.scala 137:46]
  wire [4:0] _GEN_29 = data_strb_r[0] ? 5'h8 : dc_mode_r; // @[dma.scala 131:37 dma.scala 132:33 dma.scala 34:30]
  wire [63:0] _GEN_30 = data_strb_r[0] ? data_buf_r : dc_wdata_r; // @[dma.scala 131:37 dma.scala 133:33 dma.scala 33:30]
  wire [7:0] _GEN_31 = data_strb_r[0] ? data_strb_r : _data_strb_r_T; // @[dma.scala 131:37 dma.scala 36:30 dma.scala 135:33]
  wire [63:0] _GEN_32 = data_strb_r[0] ? data_buf_r : _data_buf_r_T; // @[dma.scala 131:37 dma.scala 35:30 dma.scala 136:33]
  wire [31:0] _GEN_33 = data_strb_r[0] ? dc_addr_r : _dc_addr_r_T_13; // @[dma.scala 131:37 dma.scala 32:30 dma.scala 137:33]
  wire [4:0] _GEN_35 = _T_4 ? 5'h0 : _GEN_29; // @[dma.scala 140:62 dma.scala 141:33]
  wire [7:0] _GEN_36 = _T_4 ? _data_strb_r_T : _GEN_31; // @[dma.scala 140:62 dma.scala 142:33]
  wire [63:0] _GEN_37 = _T_4 ? _data_buf_r_T : _GEN_32; // @[dma.scala 140:62 dma.scala 143:33]
  wire [31:0] _GEN_38 = _T_4 ? _dc_addr_r_T_13 : _GEN_33; // @[dma.scala 140:62 dma.scala 144:33]
  wire [31:0] _GEN_40 = data_strb_r == 8'h0 ? _dc_addr_r_T_3 : addr_r; // @[dma.scala 117:38 dma.scala 118:24 dma.scala 39:30]
  wire [31:0] _GEN_41 = data_strb_r == 8'h0 ? _dc_addr_r_T_5 : _GEN_38; // @[dma.scala 117:38 dma.scala 119:27]
  wire  _GEN_42 = data_strb_r == 8'h0 ? _GEN_23 : bvalid_r; // @[dma.scala 117:38 dma.scala 22:30]
  wire [3:0] _GEN_44 = data_strb_r == 8'h0 ? _GEN_25 : bid_r; // @[dma.scala 117:38 dma.scala 24:30]
  wire [2:0] _GEN_45 = data_strb_r == 8'h0 ? _GEN_26 : state; // @[dma.scala 117:38 dma.scala 18:24]
  wire  _GEN_46 = data_strb_r == 8'h0 ? _GEN_27 : wready_r; // @[dma.scala 117:38 dma.scala 21:30]
  wire [7:0] _GEN_47 = data_strb_r == 8'h0 ? _GEN_28 : len_r; // @[dma.scala 117:38 dma.scala 41:30]
  wire [4:0] _GEN_48 = data_strb_r == 8'h0 ? dc_mode_r : _GEN_35; // @[dma.scala 117:38 dma.scala 34:30]
  wire [63:0] _GEN_49 = data_strb_r == 8'h0 ? dc_wdata_r : _GEN_30; // @[dma.scala 117:38 dma.scala 33:30]
  wire [7:0] _GEN_50 = data_strb_r == 8'h0 ? data_strb_r : _GEN_36; // @[dma.scala 117:38 dma.scala 36:30]
  wire [63:0] _GEN_51 = data_strb_r == 8'h0 ? data_buf_r : _GEN_37; // @[dma.scala 117:38 dma.scala 35:30]
  wire  _T_16 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_53 = io_dmaAxi_bready & bvalid_r ? 3'h0 : state; // @[dma.scala 150:47 dma.scala 151:23 dma.scala 18:24]
  wire [2:0] _GEN_55 = _T_16 ? _GEN_53 : state; // @[Conditional.scala 39:67 dma.scala 18:24]
  wire [31:0] _GEN_57 = _T_10 ? _GEN_40 : addr_r; // @[Conditional.scala 39:67 dma.scala 39:30]
  wire [31:0] _GEN_58 = _T_10 ? _GEN_41 : dc_addr_r; // @[Conditional.scala 39:67 dma.scala 32:30]
  wire  _GEN_59 = _T_10 ? _GEN_42 : bvalid_r; // @[Conditional.scala 39:67 dma.scala 22:30]
  wire [3:0] _GEN_61 = _T_10 ? _GEN_44 : bid_r; // @[Conditional.scala 39:67 dma.scala 24:30]
  wire [2:0] _GEN_62 = _T_10 ? _GEN_45 : _GEN_55; // @[Conditional.scala 39:67]
  wire  _GEN_63 = _T_10 ? _GEN_46 : wready_r; // @[Conditional.scala 39:67 dma.scala 21:30]
  wire [7:0] _GEN_64 = _T_10 ? _GEN_47 : len_r; // @[Conditional.scala 39:67 dma.scala 41:30]
  wire [4:0] _GEN_65 = _T_10 ? _GEN_48 : dc_mode_r; // @[Conditional.scala 39:67 dma.scala 34:30]
  wire [63:0] _GEN_66 = _T_10 ? _GEN_49 : dc_wdata_r; // @[Conditional.scala 39:67 dma.scala 33:30]
  wire [7:0] _GEN_67 = _T_10 ? _GEN_50 : data_strb_r; // @[Conditional.scala 39:67 dma.scala 36:30]
  wire [63:0] _GEN_68 = _T_10 ? _GEN_51 : data_buf_r; // @[Conditional.scala 39:67 dma.scala 35:30]
  wire  _GEN_70 = _T_8 ? _GEN_18 : _GEN_63; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_71 = _T_8 ? _GEN_19 : _GEN_68; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_72 = _T_8 ? _GEN_20 : _GEN_67; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_74 = _T_8 ? _GEN_22 : _GEN_62; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_75 = _T_8 ? addr_r : _GEN_57; // @[Conditional.scala 39:67 dma.scala 39:30]
  wire [31:0] _GEN_76 = _T_8 ? dc_addr_r : _GEN_58; // @[Conditional.scala 39:67 dma.scala 32:30]
  wire  _GEN_77 = _T_8 ? bvalid_r : _GEN_59; // @[Conditional.scala 39:67 dma.scala 22:30]
  wire [3:0] _GEN_79 = _T_8 ? bid_r : _GEN_61; // @[Conditional.scala 39:67 dma.scala 24:30]
  wire [7:0] _GEN_80 = _T_8 ? len_r : _GEN_64; // @[Conditional.scala 39:67 dma.scala 41:30]
  wire [4:0] _GEN_81 = _T_8 ? dc_mode_r : _GEN_65; // @[Conditional.scala 39:67 dma.scala 34:30]
  wire [63:0] _GEN_82 = _T_8 ? dc_wdata_r : _GEN_66; // @[Conditional.scala 39:67 dma.scala 33:30]
  wire  _GEN_83 = _T_7 ? 1'h0 : awready_r; // @[Conditional.scala 39:67 dma.scala 97:25 dma.scala 20:30]
  wire [31:0] _GEN_84 = _T_7 ? io_dmaAxi_awaddr : _GEN_75; // @[Conditional.scala 39:67 dma.scala 98:25]
  wire [31:0] _GEN_85 = _T_7 ? _dc_addr_r_T_7 : _GEN_76; // @[Conditional.scala 39:67 dma.scala 99:25]
  wire [3:0] _GEN_86 = _T_7 ? io_dmaAxi_awid : id_r; // @[Conditional.scala 39:67 dma.scala 100:25 dma.scala 40:30]
  wire [7:0] _GEN_87 = _T_7 ? io_dmaAxi_awlen : _GEN_80; // @[Conditional.scala 39:67 dma.scala 101:25]
  wire [7:0] _GEN_88 = _T_7 ? _size_r_T_1 : size_r; // @[Conditional.scala 39:67 dma.scala 102:25 dma.scala 42:30]
  wire  _GEN_90 = _T_7 | _GEN_70; // @[Conditional.scala 39:67 dma.scala 104:25]
  wire [2:0] _GEN_91 = _T_7 ? 3'h4 : _GEN_74; // @[Conditional.scala 39:67 dma.scala 105:25]
  wire [63:0] _GEN_92 = _T_7 ? data_buf_r : _GEN_71; // @[Conditional.scala 39:67 dma.scala 35:30]
  wire [7:0] _GEN_93 = _T_7 ? data_strb_r : _GEN_72; // @[Conditional.scala 39:67 dma.scala 36:30]
  wire  _GEN_95 = _T_7 ? bvalid_r : _GEN_77; // @[Conditional.scala 39:67 dma.scala 22:30]
  wire [3:0] _GEN_97 = _T_7 ? bid_r : _GEN_79; // @[Conditional.scala 39:67 dma.scala 24:30]
  wire [4:0] _GEN_98 = _T_7 ? dc_mode_r : _GEN_81; // @[Conditional.scala 39:67 dma.scala 34:30]
  wire [63:0] _GEN_99 = _T_7 ? dc_wdata_r : _GEN_82; // @[Conditional.scala 39:67 dma.scala 33:30]
  wire [63:0] _GEN_100 = _T_5 ? data_buf_r : rdata_r; // @[Conditional.scala 39:67 dma.scala 78:21 dma.scala 28:30]
  wire  _GEN_101 = _T_5 ? _GEN_12 : rvalid_r; // @[Conditional.scala 39:67 dma.scala 26:30]
  wire  _GEN_102 = _T_5 ? len_r == 8'h0 : rlast_r; // @[Conditional.scala 39:67 dma.scala 80:21 dma.scala 29:30]
  wire [3:0] _GEN_103 = _T_5 ? id_r : rid_r; // @[Conditional.scala 39:67 dma.scala 81:21 dma.scala 30:30]
  wire [2:0] _GEN_105 = _T_5 ? _GEN_13 : _GEN_91; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_106 = _T_5 ? _GEN_14 : _GEN_87; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_107 = _T_5 ? _GEN_15 : _GEN_85; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_108 = _T_5 ? _GEN_16 : _GEN_84; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_109 = _T_5 ? _GEN_17 : _GEN_98; // @[Conditional.scala 39:67]
  wire  _GEN_110 = _T_5 ? awready_r : _GEN_83; // @[Conditional.scala 39:67 dma.scala 20:30]
  wire [3:0] _GEN_111 = _T_5 ? id_r : _GEN_86; // @[Conditional.scala 39:67 dma.scala 40:30]
  wire [7:0] _GEN_112 = _T_5 ? size_r : _GEN_88; // @[Conditional.scala 39:67 dma.scala 42:30]
  wire  _GEN_114 = _T_5 ? wready_r : _GEN_90; // @[Conditional.scala 39:67 dma.scala 21:30]
  wire [63:0] _GEN_115 = _T_5 ? data_buf_r : _GEN_92; // @[Conditional.scala 39:67 dma.scala 35:30]
  wire [7:0] _GEN_116 = _T_5 ? data_strb_r : _GEN_93; // @[Conditional.scala 39:67 dma.scala 36:30]
  wire  _GEN_118 = _T_5 ? bvalid_r : _GEN_95; // @[Conditional.scala 39:67 dma.scala 22:30]
  wire [3:0] _GEN_120 = _T_5 ? bid_r : _GEN_97; // @[Conditional.scala 39:67 dma.scala 24:30]
  wire [63:0] _GEN_121 = _T_5 ? dc_wdata_r : _GEN_99; // @[Conditional.scala 39:67 dma.scala 33:30]
  assign io_dmaAxi_awready = awready_r; // @[dma.scala 156:25]
  assign io_dmaAxi_wready = wready_r; // @[dma.scala 157:25]
  assign io_dmaAxi_bvalid = bvalid_r; // @[dma.scala 158:25]
  assign io_dmaAxi_bid = bid_r; // @[dma.scala 160:25]
  assign io_dmaAxi_arready = arready_r; // @[dma.scala 161:25]
  assign io_dmaAxi_rvalid = rvalid_r; // @[dma.scala 162:25]
  assign io_dmaAxi_rdata = rdata_r; // @[dma.scala 164:25]
  assign io_dmaAxi_rlast = rlast_r; // @[dma.scala 165:25]
  assign io_dmaAxi_rid = rid_r; // @[dma.scala 166:25]
  assign io_dcRW_addr = dc_addr_r; // @[dma.scala 168:21]
  assign io_dcRW_wdata = dc_wdata_r; // @[dma.scala 169:21]
  assign io_dcRW_dc_mode = dc_mode_r; // @[dma.scala 170:21]
  always @(posedge clock) begin
    if (reset) begin // @[dma.scala 18:24]
      state <= 3'h0; // @[dma.scala 18:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_dmaAxi_awvalid) begin // @[dma.scala 52:36]
        state <= 3'h3; // @[dma.scala 53:29]
      end else if (io_dmaAxi_arvalid) begin // @[dma.scala 48:36]
        state <= 3'h1; // @[dma.scala 49:29]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      state <= 3'h6; // @[dma.scala 64:25]
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      state <= _GEN_6;
    end else begin
      state <= _GEN_105;
    end
    if (reset) begin // @[dma.scala 20:30]
      awready_r <= 1'h0; // @[dma.scala 20:30]
    end else if (_T) begin // @[Conditional.scala 40:58]
      awready_r <= _GEN_3;
    end else if (!(_T_1)) begin // @[Conditional.scala 39:67]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        awready_r <= _GEN_110;
      end
    end
    if (reset) begin // @[dma.scala 21:30]
      wready_r <= 1'h0; // @[dma.scala 21:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          wready_r <= _GEN_114;
        end
      end
    end
    if (reset) begin // @[dma.scala 22:30]
      bvalid_r <= 1'h0; // @[dma.scala 22:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          bvalid_r <= _GEN_118;
        end
      end
    end
    if (reset) begin // @[dma.scala 24:30]
      bid_r <= 4'h0; // @[dma.scala 24:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          bid_r <= _GEN_120;
        end
      end
    end
    if (reset) begin // @[dma.scala 25:30]
      arready_r <= 1'h0; // @[dma.scala 25:30]
    end else if (_T) begin // @[Conditional.scala 40:58]
      arready_r <= _GEN_1;
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      arready_r <= 1'h0; // @[dma.scala 58:25]
    end
    if (reset) begin // @[dma.scala 26:30]
      rvalid_r <= 1'h0; // @[dma.scala 26:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          rvalid_r <= _GEN_101;
        end
      end
    end
    if (reset) begin // @[dma.scala 28:30]
      rdata_r <= 64'h0; // @[dma.scala 28:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          rdata_r <= _GEN_100;
        end
      end
    end
    if (reset) begin // @[dma.scala 29:30]
      rlast_r <= 1'h0; // @[dma.scala 29:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          rlast_r <= _GEN_102;
        end
      end
    end
    if (reset) begin // @[dma.scala 30:30]
      rid_r <= 4'h0; // @[dma.scala 30:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          rid_r <= _GEN_103;
        end
      end
    end
    if (reset) begin // @[dma.scala 32:30]
      dc_addr_r <= 32'h0; // @[dma.scala 32:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        dc_addr_r <= _dc_addr_r_T_1; // @[dma.scala 65:25]
      end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
        dc_addr_r <= _GEN_107;
      end
    end
    if (reset) begin // @[dma.scala 33:30]
      dc_wdata_r <= 64'h0; // @[dma.scala 33:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          dc_wdata_r <= _GEN_121;
        end
      end
    end
    if (reset) begin // @[dma.scala 34:30]
      dc_mode_r <= 5'h0; // @[dma.scala 34:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        dc_mode_r <= 5'h7; // @[dma.scala 66:25]
      end else if (_T_2) begin // @[Conditional.scala 39:67]
        dc_mode_r <= _GEN_4;
      end else begin
        dc_mode_r <= _GEN_109;
      end
    end
    if (reset) begin // @[dma.scala 35:30]
      data_buf_r <= 64'h0; // @[dma.scala 35:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          data_buf_r <= _GEN_5;
        end else begin
          data_buf_r <= _GEN_115;
        end
      end
    end
    if (reset) begin // @[dma.scala 36:30]
      data_strb_r <= 8'h0; // @[dma.scala 36:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          data_strb_r <= _GEN_116;
        end
      end
    end
    if (reset) begin // @[dma.scala 39:30]
      addr_r <= 32'h0; // @[dma.scala 39:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        addr_r <= io_dmaAxi_araddr; // @[dma.scala 59:25]
      end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
        addr_r <= _GEN_108;
      end
    end
    if (reset) begin // @[dma.scala 40:30]
      id_r <= 4'h0; // @[dma.scala 40:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        id_r <= io_dmaAxi_arid; // @[dma.scala 60:25]
      end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
        id_r <= _GEN_111;
      end
    end
    if (reset) begin // @[dma.scala 41:30]
      len_r <= 8'h0; // @[dma.scala 41:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        len_r <= io_dmaAxi_arlen; // @[dma.scala 61:25]
      end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
        len_r <= _GEN_106;
      end
    end
    if (reset) begin // @[dma.scala 42:30]
      size_r <= 8'h0; // @[dma.scala 42:30]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        size_r <= _size_r_T; // @[dma.scala 62:25]
      end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
        size_r <= _GEN_112;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  awready_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wready_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bvalid_r = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bid_r = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  arready_r = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  rvalid_r = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  rdata_r = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  rlast_r = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  rid_r = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  dc_addr_r = _RAND_10[31:0];
  _RAND_11 = {2{`RANDOM}};
  dc_wdata_r = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  dc_mode_r = _RAND_12[4:0];
  _RAND_13 = {2{`RANDOM}};
  data_buf_r = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  data_strb_r = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  addr_r = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  id_r = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  len_r = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  size_r = _RAND_18[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_000000(
  input          clock,
  input          reset,
  input          io_master_awready,
  output         io_master_awvalid,
  output [31:0]  io_master_awaddr,
  output [3:0]   io_master_awid,
  output [7:0]   io_master_awlen,
  output [2:0]   io_master_awsize,
  output [1:0]   io_master_awburst,
  input          io_master_wready,
  output         io_master_wvalid,
  output [63:0]  io_master_wdata,
  output [7:0]   io_master_wstrb,
  output         io_master_wlast,
  output         io_master_bready,
  input          io_master_bvalid,
  input  [1:0]   io_master_bresp,
  input  [3:0]   io_master_bid,
  input          io_master_arready,
  output         io_master_arvalid,
  output [31:0]  io_master_araddr,
  output [3:0]   io_master_arid,
  output [7:0]   io_master_arlen,
  output [2:0]   io_master_arsize,
  output [1:0]   io_master_arburst,
  output         io_master_rready,
  input          io_master_rvalid,
  input  [1:0]   io_master_rresp,
  input  [63:0]  io_master_rdata,
  input          io_master_rlast,
  input  [3:0]   io_master_rid,
  output         io_slave_awready,
  input          io_slave_awvalid,
  input  [31:0]  io_slave_awaddr,
  input  [3:0]   io_slave_awid,
  input  [7:0]   io_slave_awlen,
  input  [2:0]   io_slave_awsize,
  input  [1:0]   io_slave_awburst,
  output         io_slave_wready,
  input          io_slave_wvalid,
  input  [63:0]  io_slave_wdata,
  input  [7:0]   io_slave_wstrb,
  input          io_slave_wlast,
  input          io_slave_bready,
  output         io_slave_bvalid,
  output [1:0]   io_slave_bresp,
  output [3:0]   io_slave_bid,
  output         io_slave_arready,
  input          io_slave_arvalid,
  input  [31:0]  io_slave_araddr,
  input  [3:0]   io_slave_arid,
  input  [7:0]   io_slave_arlen,
  input  [2:0]   io_slave_arsize,
  input  [1:0]   io_slave_arburst,
  input          io_slave_rready,
  output         io_slave_rvalid,
  output [1:0]   io_slave_rresp,
  output [63:0]  io_slave_rdata,
  output         io_slave_rlast,
  output [3:0]   io_slave_rid,
  output [5:0]   io_sram0_addr,
  output         io_sram0_cen,
  output         io_sram0_wen,
  output [127:0] io_sram0_wmask,
  output [127:0] io_sram0_wdata,
  input  [127:0] io_sram0_rdata,
  output [5:0]   io_sram1_addr,
  output         io_sram1_cen,
  output         io_sram1_wen,
  output [127:0] io_sram1_wmask,
  output [127:0] io_sram1_wdata,
  input  [127:0] io_sram1_rdata,
  output [5:0]   io_sram2_addr,
  output         io_sram2_cen,
  output         io_sram2_wen,
  output [127:0] io_sram2_wmask,
  output [127:0] io_sram2_wdata,
  input  [127:0] io_sram2_rdata,
  output [5:0]   io_sram3_addr,
  output         io_sram3_cen,
  output         io_sram3_wen,
  output [127:0] io_sram3_wmask,
  output [127:0] io_sram3_wdata,
  input  [127:0] io_sram3_rdata,
  output [5:0]   io_sram4_addr,
  output         io_sram4_cen,
  output         io_sram4_wen,
  output [127:0] io_sram4_wmask,
  output [127:0] io_sram4_wdata,
  input  [127:0] io_sram4_rdata,
  output [5:0]   io_sram5_addr,
  output         io_sram5_cen,
  output         io_sram5_wen,
  output [127:0] io_sram5_wmask,
  output [127:0] io_sram5_wdata,
  input  [127:0] io_sram5_rdata,
  output [5:0]   io_sram6_addr,
  output         io_sram6_cen,
  output         io_sram6_wen,
  output [127:0] io_sram6_wmask,
  output [127:0] io_sram6_wdata,
  input  [127:0] io_sram6_rdata,
  output [5:0]   io_sram7_addr,
  output         io_sram7_cen,
  output         io_sram7_wen,
  output [127:0] io_sram7_wmask,
  output [127:0] io_sram7_wdata,
  input  [127:0] io_sram7_rdata,
  input          io_interrupt
);
  wire  fetch_clock; // @[cpu.scala 71:29]
  wire  fetch_reset; // @[cpu.scala 71:29]
  wire [31:0] fetch_io_instRead_addr; // @[cpu.scala 71:29]
  wire [63:0] fetch_io_instRead_inst; // @[cpu.scala 71:29]
  wire  fetch_io_instRead_arvalid; // @[cpu.scala 71:29]
  wire  fetch_io_instRead_rvalid; // @[cpu.scala 71:29]
  wire [63:0] fetch_io_va2pa_vaddr; // @[cpu.scala 71:29]
  wire  fetch_io_va2pa_vvalid; // @[cpu.scala 71:29]
  wire [31:0] fetch_io_va2pa_paddr; // @[cpu.scala 71:29]
  wire  fetch_io_va2pa_pvalid; // @[cpu.scala 71:29]
  wire [63:0] fetch_io_va2pa_tlb_excep_cause; // @[cpu.scala 71:29]
  wire [63:0] fetch_io_va2pa_tlb_excep_tval; // @[cpu.scala 71:29]
  wire  fetch_io_va2pa_tlb_excep_en; // @[cpu.scala 71:29]
  wire [63:0] fetch_io_reg2if_seq_pc; // @[cpu.scala 71:29]
  wire  fetch_io_reg2if_valid; // @[cpu.scala 71:29]
  wire [63:0] fetch_io_wb2if_seq_pc; // @[cpu.scala 71:29]
  wire  fetch_io_wb2if_valid; // @[cpu.scala 71:29]
  wire  fetch_io_recov; // @[cpu.scala 71:29]
  wire  fetch_io_intr_in_en; // @[cpu.scala 71:29]
  wire [63:0] fetch_io_intr_in_cause; // @[cpu.scala 71:29]
  wire [63:0] fetch_io_branchFail_seq_pc; // @[cpu.scala 71:29]
  wire  fetch_io_branchFail_valid; // @[cpu.scala 71:29]
  wire [31:0] fetch_io_if2id_inst; // @[cpu.scala 71:29]
  wire [63:0] fetch_io_if2id_pc; // @[cpu.scala 71:29]
  wire [63:0] fetch_io_if2id_excep_cause; // @[cpu.scala 71:29]
  wire [63:0] fetch_io_if2id_excep_tval; // @[cpu.scala 71:29]
  wire  fetch_io_if2id_excep_en; // @[cpu.scala 71:29]
  wire [63:0] fetch_io_if2id_excep_pc; // @[cpu.scala 71:29]
  wire  fetch_io_if2id_drop; // @[cpu.scala 71:29]
  wire  fetch_io_if2id_stall; // @[cpu.scala 71:29]
  wire  fetch_io_if2id_recov; // @[cpu.scala 71:29]
  wire  fetch_io_if2id_valid; // @[cpu.scala 71:29]
  wire  fetch_io_if2id_ready; // @[cpu.scala 71:29]
  wire  decode_clock; // @[cpu.scala 72:29]
  wire  decode_reset; // @[cpu.scala 72:29]
  wire [31:0] decode_io_if2id_inst; // @[cpu.scala 72:29]
  wire [63:0] decode_io_if2id_pc; // @[cpu.scala 72:29]
  wire [63:0] decode_io_if2id_excep_cause; // @[cpu.scala 72:29]
  wire [63:0] decode_io_if2id_excep_tval; // @[cpu.scala 72:29]
  wire  decode_io_if2id_excep_en; // @[cpu.scala 72:29]
  wire [63:0] decode_io_if2id_excep_pc; // @[cpu.scala 72:29]
  wire  decode_io_if2id_drop; // @[cpu.scala 72:29]
  wire  decode_io_if2id_stall; // @[cpu.scala 72:29]
  wire  decode_io_if2id_recov; // @[cpu.scala 72:29]
  wire  decode_io_if2id_valid; // @[cpu.scala 72:29]
  wire  decode_io_if2id_ready; // @[cpu.scala 72:29]
  wire [31:0] decode_io_id2df_inst; // @[cpu.scala 72:29]
  wire [63:0] decode_io_id2df_pc; // @[cpu.scala 72:29]
  wire [63:0] decode_io_id2df_excep_cause; // @[cpu.scala 72:29]
  wire [63:0] decode_io_id2df_excep_tval; // @[cpu.scala 72:29]
  wire  decode_io_id2df_excep_en; // @[cpu.scala 72:29]
  wire [63:0] decode_io_id2df_excep_pc; // @[cpu.scala 72:29]
  wire [1:0] decode_io_id2df_excep_etype; // @[cpu.scala 72:29]
  wire [4:0] decode_io_id2df_ctrl_aluOp; // @[cpu.scala 72:29]
  wire  decode_io_id2df_ctrl_aluWidth; // @[cpu.scala 72:29]
  wire [4:0] decode_io_id2df_ctrl_dcMode; // @[cpu.scala 72:29]
  wire  decode_io_id2df_ctrl_writeRegEn; // @[cpu.scala 72:29]
  wire  decode_io_id2df_ctrl_writeCSREn; // @[cpu.scala 72:29]
  wire [2:0] decode_io_id2df_ctrl_brType; // @[cpu.scala 72:29]
  wire [4:0] decode_io_id2df_rs1; // @[cpu.scala 72:29]
  wire  decode_io_id2df_rrs1; // @[cpu.scala 72:29]
  wire [63:0] decode_io_id2df_rs1_d; // @[cpu.scala 72:29]
  wire [11:0] decode_io_id2df_rs2; // @[cpu.scala 72:29]
  wire  decode_io_id2df_rrs2; // @[cpu.scala 72:29]
  wire [63:0] decode_io_id2df_rs2_d; // @[cpu.scala 72:29]
  wire [4:0] decode_io_id2df_dst; // @[cpu.scala 72:29]
  wire [63:0] decode_io_id2df_dst_d; // @[cpu.scala 72:29]
  wire [1:0] decode_io_id2df_jmp_type; // @[cpu.scala 72:29]
  wire [1:0] decode_io_id2df_special; // @[cpu.scala 72:29]
  wire [5:0] decode_io_id2df_swap; // @[cpu.scala 72:29]
  wire [1:0] decode_io_id2df_indi; // @[cpu.scala 72:29]
  wire  decode_io_id2df_drop; // @[cpu.scala 72:29]
  wire  decode_io_id2df_stall; // @[cpu.scala 72:29]
  wire  decode_io_id2df_recov; // @[cpu.scala 72:29]
  wire  decode_io_id2df_valid; // @[cpu.scala 72:29]
  wire  decode_io_id2df_ready; // @[cpu.scala 72:29]
  wire [1:0] decode_io_idState_priv; // @[cpu.scala 72:29]
  wire  forwading_clock; // @[cpu.scala 73:29]
  wire  forwading_reset; // @[cpu.scala 73:29]
  wire [31:0] forwading_io_id2df_inst; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_id2df_pc; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_id2df_excep_cause; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_id2df_excep_tval; // @[cpu.scala 73:29]
  wire  forwading_io_id2df_excep_en; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_id2df_excep_pc; // @[cpu.scala 73:29]
  wire [1:0] forwading_io_id2df_excep_etype; // @[cpu.scala 73:29]
  wire [4:0] forwading_io_id2df_ctrl_aluOp; // @[cpu.scala 73:29]
  wire  forwading_io_id2df_ctrl_aluWidth; // @[cpu.scala 73:29]
  wire [4:0] forwading_io_id2df_ctrl_dcMode; // @[cpu.scala 73:29]
  wire  forwading_io_id2df_ctrl_writeRegEn; // @[cpu.scala 73:29]
  wire  forwading_io_id2df_ctrl_writeCSREn; // @[cpu.scala 73:29]
  wire [2:0] forwading_io_id2df_ctrl_brType; // @[cpu.scala 73:29]
  wire [4:0] forwading_io_id2df_rs1; // @[cpu.scala 73:29]
  wire  forwading_io_id2df_rrs1; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_id2df_rs1_d; // @[cpu.scala 73:29]
  wire [11:0] forwading_io_id2df_rs2; // @[cpu.scala 73:29]
  wire  forwading_io_id2df_rrs2; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_id2df_rs2_d; // @[cpu.scala 73:29]
  wire [4:0] forwading_io_id2df_dst; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_id2df_dst_d; // @[cpu.scala 73:29]
  wire [1:0] forwading_io_id2df_jmp_type; // @[cpu.scala 73:29]
  wire [1:0] forwading_io_id2df_special; // @[cpu.scala 73:29]
  wire [5:0] forwading_io_id2df_swap; // @[cpu.scala 73:29]
  wire [1:0] forwading_io_id2df_indi; // @[cpu.scala 73:29]
  wire  forwading_io_id2df_drop; // @[cpu.scala 73:29]
  wire  forwading_io_id2df_stall; // @[cpu.scala 73:29]
  wire  forwading_io_id2df_recov; // @[cpu.scala 73:29]
  wire  forwading_io_id2df_valid; // @[cpu.scala 73:29]
  wire  forwading_io_id2df_ready; // @[cpu.scala 73:29]
  wire [31:0] forwading_io_df2rr_inst; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_df2rr_pc; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_df2rr_excep_cause; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_df2rr_excep_tval; // @[cpu.scala 73:29]
  wire  forwading_io_df2rr_excep_en; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_df2rr_excep_pc; // @[cpu.scala 73:29]
  wire [1:0] forwading_io_df2rr_excep_etype; // @[cpu.scala 73:29]
  wire [4:0] forwading_io_df2rr_ctrl_aluOp; // @[cpu.scala 73:29]
  wire  forwading_io_df2rr_ctrl_aluWidth; // @[cpu.scala 73:29]
  wire [4:0] forwading_io_df2rr_ctrl_dcMode; // @[cpu.scala 73:29]
  wire  forwading_io_df2rr_ctrl_writeRegEn; // @[cpu.scala 73:29]
  wire  forwading_io_df2rr_ctrl_writeCSREn; // @[cpu.scala 73:29]
  wire [2:0] forwading_io_df2rr_ctrl_brType; // @[cpu.scala 73:29]
  wire [4:0] forwading_io_df2rr_rs1; // @[cpu.scala 73:29]
  wire  forwading_io_df2rr_rrs1; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_df2rr_rs1_d; // @[cpu.scala 73:29]
  wire [11:0] forwading_io_df2rr_rs2; // @[cpu.scala 73:29]
  wire  forwading_io_df2rr_rrs2; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_df2rr_rs2_d; // @[cpu.scala 73:29]
  wire [4:0] forwading_io_df2rr_dst; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_df2rr_dst_d; // @[cpu.scala 73:29]
  wire [1:0] forwading_io_df2rr_jmp_type; // @[cpu.scala 73:29]
  wire [1:0] forwading_io_df2rr_special; // @[cpu.scala 73:29]
  wire [5:0] forwading_io_df2rr_swap; // @[cpu.scala 73:29]
  wire [1:0] forwading_io_df2rr_indi; // @[cpu.scala 73:29]
  wire  forwading_io_df2rr_drop; // @[cpu.scala 73:29]
  wire  forwading_io_df2rr_stall; // @[cpu.scala 73:29]
  wire  forwading_io_df2rr_recov; // @[cpu.scala 73:29]
  wire  forwading_io_df2rr_valid; // @[cpu.scala 73:29]
  wire  forwading_io_df2rr_ready; // @[cpu.scala 73:29]
  wire [4:0] forwading_io_d_rr_id; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_d_rr_data; // @[cpu.scala 73:29]
  wire [1:0] forwading_io_d_rr_state; // @[cpu.scala 73:29]
  wire [4:0] forwading_io_d_ex_id; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_d_ex_data; // @[cpu.scala 73:29]
  wire [1:0] forwading_io_d_ex_state; // @[cpu.scala 73:29]
  wire [4:0] forwading_io_d_mem1_id; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_d_mem1_data; // @[cpu.scala 73:29]
  wire [1:0] forwading_io_d_mem1_state; // @[cpu.scala 73:29]
  wire [4:0] forwading_io_d_mem2_id; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_d_mem2_data; // @[cpu.scala 73:29]
  wire [1:0] forwading_io_d_mem2_state; // @[cpu.scala 73:29]
  wire [4:0] forwading_io_d_mem3_id; // @[cpu.scala 73:29]
  wire [63:0] forwading_io_d_mem3_data; // @[cpu.scala 73:29]
  wire [1:0] forwading_io_d_mem3_state; // @[cpu.scala 73:29]
  wire  readregs_clock; // @[cpu.scala 74:29]
  wire  readregs_reset; // @[cpu.scala 74:29]
  wire [31:0] readregs_io_df2rr_inst; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_df2rr_pc; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_df2rr_excep_cause; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_df2rr_excep_tval; // @[cpu.scala 74:29]
  wire  readregs_io_df2rr_excep_en; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_df2rr_excep_pc; // @[cpu.scala 74:29]
  wire [1:0] readregs_io_df2rr_excep_etype; // @[cpu.scala 74:29]
  wire [4:0] readregs_io_df2rr_ctrl_aluOp; // @[cpu.scala 74:29]
  wire  readregs_io_df2rr_ctrl_aluWidth; // @[cpu.scala 74:29]
  wire [4:0] readregs_io_df2rr_ctrl_dcMode; // @[cpu.scala 74:29]
  wire  readregs_io_df2rr_ctrl_writeRegEn; // @[cpu.scala 74:29]
  wire  readregs_io_df2rr_ctrl_writeCSREn; // @[cpu.scala 74:29]
  wire [2:0] readregs_io_df2rr_ctrl_brType; // @[cpu.scala 74:29]
  wire [4:0] readregs_io_df2rr_rs1; // @[cpu.scala 74:29]
  wire  readregs_io_df2rr_rrs1; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_df2rr_rs1_d; // @[cpu.scala 74:29]
  wire [11:0] readregs_io_df2rr_rs2; // @[cpu.scala 74:29]
  wire  readregs_io_df2rr_rrs2; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_df2rr_rs2_d; // @[cpu.scala 74:29]
  wire [4:0] readregs_io_df2rr_dst; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_df2rr_dst_d; // @[cpu.scala 74:29]
  wire [1:0] readregs_io_df2rr_jmp_type; // @[cpu.scala 74:29]
  wire [1:0] readregs_io_df2rr_special; // @[cpu.scala 74:29]
  wire [5:0] readregs_io_df2rr_swap; // @[cpu.scala 74:29]
  wire [1:0] readregs_io_df2rr_indi; // @[cpu.scala 74:29]
  wire  readregs_io_df2rr_drop; // @[cpu.scala 74:29]
  wire  readregs_io_df2rr_stall; // @[cpu.scala 74:29]
  wire  readregs_io_df2rr_recov; // @[cpu.scala 74:29]
  wire  readregs_io_df2rr_valid; // @[cpu.scala 74:29]
  wire  readregs_io_df2rr_ready; // @[cpu.scala 74:29]
  wire [31:0] readregs_io_rr2ex_inst; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_rr2ex_pc; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_rr2ex_excep_cause; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_rr2ex_excep_tval; // @[cpu.scala 74:29]
  wire  readregs_io_rr2ex_excep_en; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_rr2ex_excep_pc; // @[cpu.scala 74:29]
  wire [1:0] readregs_io_rr2ex_excep_etype; // @[cpu.scala 74:29]
  wire [4:0] readregs_io_rr2ex_ctrl_aluOp; // @[cpu.scala 74:29]
  wire  readregs_io_rr2ex_ctrl_aluWidth; // @[cpu.scala 74:29]
  wire [4:0] readregs_io_rr2ex_ctrl_dcMode; // @[cpu.scala 74:29]
  wire  readregs_io_rr2ex_ctrl_writeRegEn; // @[cpu.scala 74:29]
  wire  readregs_io_rr2ex_ctrl_writeCSREn; // @[cpu.scala 74:29]
  wire [2:0] readregs_io_rr2ex_ctrl_brType; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_rr2ex_rs1_d; // @[cpu.scala 74:29]
  wire [11:0] readregs_io_rr2ex_rs2; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_rr2ex_rs2_d; // @[cpu.scala 74:29]
  wire [4:0] readregs_io_rr2ex_dst; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_rr2ex_dst_d; // @[cpu.scala 74:29]
  wire [11:0] readregs_io_rr2ex_rcsr_id; // @[cpu.scala 74:29]
  wire [1:0] readregs_io_rr2ex_jmp_type; // @[cpu.scala 74:29]
  wire [1:0] readregs_io_rr2ex_special; // @[cpu.scala 74:29]
  wire [1:0] readregs_io_rr2ex_indi; // @[cpu.scala 74:29]
  wire  readregs_io_rr2ex_drop; // @[cpu.scala 74:29]
  wire  readregs_io_rr2ex_stall; // @[cpu.scala 74:29]
  wire  readregs_io_rr2ex_recov; // @[cpu.scala 74:29]
  wire  readregs_io_rr2ex_valid; // @[cpu.scala 74:29]
  wire  readregs_io_rr2ex_ready; // @[cpu.scala 74:29]
  wire [4:0] readregs_io_rs1Read_id; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_rs1Read_data; // @[cpu.scala 74:29]
  wire [4:0] readregs_io_rs2Read_id; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_rs2Read_data; // @[cpu.scala 74:29]
  wire [11:0] readregs_io_csrRead_id; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_csrRead_data; // @[cpu.scala 74:29]
  wire  readregs_io_csrRead_is_err; // @[cpu.scala 74:29]
  wire [4:0] readregs_io_d_rr_id; // @[cpu.scala 74:29]
  wire [63:0] readregs_io_d_rr_data; // @[cpu.scala 74:29]
  wire [1:0] readregs_io_d_rr_state; // @[cpu.scala 74:29]
  wire  execute_clock; // @[cpu.scala 75:29]
  wire  execute_reset; // @[cpu.scala 75:29]
  wire [31:0] execute_io_rr2ex_inst; // @[cpu.scala 75:29]
  wire [63:0] execute_io_rr2ex_pc; // @[cpu.scala 75:29]
  wire [63:0] execute_io_rr2ex_excep_cause; // @[cpu.scala 75:29]
  wire [63:0] execute_io_rr2ex_excep_tval; // @[cpu.scala 75:29]
  wire  execute_io_rr2ex_excep_en; // @[cpu.scala 75:29]
  wire [63:0] execute_io_rr2ex_excep_pc; // @[cpu.scala 75:29]
  wire [1:0] execute_io_rr2ex_excep_etype; // @[cpu.scala 75:29]
  wire [4:0] execute_io_rr2ex_ctrl_aluOp; // @[cpu.scala 75:29]
  wire  execute_io_rr2ex_ctrl_aluWidth; // @[cpu.scala 75:29]
  wire [4:0] execute_io_rr2ex_ctrl_dcMode; // @[cpu.scala 75:29]
  wire  execute_io_rr2ex_ctrl_writeRegEn; // @[cpu.scala 75:29]
  wire  execute_io_rr2ex_ctrl_writeCSREn; // @[cpu.scala 75:29]
  wire [2:0] execute_io_rr2ex_ctrl_brType; // @[cpu.scala 75:29]
  wire [63:0] execute_io_rr2ex_rs1_d; // @[cpu.scala 75:29]
  wire [11:0] execute_io_rr2ex_rs2; // @[cpu.scala 75:29]
  wire [63:0] execute_io_rr2ex_rs2_d; // @[cpu.scala 75:29]
  wire [4:0] execute_io_rr2ex_dst; // @[cpu.scala 75:29]
  wire [63:0] execute_io_rr2ex_dst_d; // @[cpu.scala 75:29]
  wire [11:0] execute_io_rr2ex_rcsr_id; // @[cpu.scala 75:29]
  wire [1:0] execute_io_rr2ex_jmp_type; // @[cpu.scala 75:29]
  wire [1:0] execute_io_rr2ex_special; // @[cpu.scala 75:29]
  wire [1:0] execute_io_rr2ex_indi; // @[cpu.scala 75:29]
  wire  execute_io_rr2ex_drop; // @[cpu.scala 75:29]
  wire  execute_io_rr2ex_stall; // @[cpu.scala 75:29]
  wire  execute_io_rr2ex_recov; // @[cpu.scala 75:29]
  wire  execute_io_rr2ex_valid; // @[cpu.scala 75:29]
  wire  execute_io_rr2ex_ready; // @[cpu.scala 75:29]
  wire [31:0] execute_io_ex2mem_inst; // @[cpu.scala 75:29]
  wire [63:0] execute_io_ex2mem_pc; // @[cpu.scala 75:29]
  wire [63:0] execute_io_ex2mem_excep_cause; // @[cpu.scala 75:29]
  wire [63:0] execute_io_ex2mem_excep_tval; // @[cpu.scala 75:29]
  wire  execute_io_ex2mem_excep_en; // @[cpu.scala 75:29]
  wire [63:0] execute_io_ex2mem_excep_pc; // @[cpu.scala 75:29]
  wire [1:0] execute_io_ex2mem_excep_etype; // @[cpu.scala 75:29]
  wire [4:0] execute_io_ex2mem_ctrl_dcMode; // @[cpu.scala 75:29]
  wire  execute_io_ex2mem_ctrl_writeRegEn; // @[cpu.scala 75:29]
  wire  execute_io_ex2mem_ctrl_writeCSREn; // @[cpu.scala 75:29]
  wire [63:0] execute_io_ex2mem_mem_addr; // @[cpu.scala 75:29]
  wire [63:0] execute_io_ex2mem_mem_data; // @[cpu.scala 75:29]
  wire [11:0] execute_io_ex2mem_csr_id; // @[cpu.scala 75:29]
  wire [63:0] execute_io_ex2mem_csr_d; // @[cpu.scala 75:29]
  wire [4:0] execute_io_ex2mem_dst; // @[cpu.scala 75:29]
  wire [63:0] execute_io_ex2mem_dst_d; // @[cpu.scala 75:29]
  wire [11:0] execute_io_ex2mem_rcsr_id; // @[cpu.scala 75:29]
  wire [1:0] execute_io_ex2mem_special; // @[cpu.scala 75:29]
  wire [1:0] execute_io_ex2mem_indi; // @[cpu.scala 75:29]
  wire  execute_io_ex2mem_drop; // @[cpu.scala 75:29]
  wire  execute_io_ex2mem_stall; // @[cpu.scala 75:29]
  wire  execute_io_ex2mem_recov; // @[cpu.scala 75:29]
  wire  execute_io_ex2mem_valid; // @[cpu.scala 75:29]
  wire  execute_io_ex2mem_ready; // @[cpu.scala 75:29]
  wire [4:0] execute_io_d_ex_id; // @[cpu.scala 75:29]
  wire [63:0] execute_io_d_ex_data; // @[cpu.scala 75:29]
  wire [1:0] execute_io_d_ex_state; // @[cpu.scala 75:29]
  wire [63:0] execute_io_ex2if_seq_pc; // @[cpu.scala 75:29]
  wire  execute_io_ex2if_valid; // @[cpu.scala 75:29]
  wire [63:0] execute_io_updateNextPc_seq_pc; // @[cpu.scala 75:29]
  wire  execute_io_updateNextPc_valid; // @[cpu.scala 75:29]
  wire  memory_clock; // @[cpu.scala 76:29]
  wire  memory_reset; // @[cpu.scala 76:29]
  wire [31:0] memory_io_ex2mem_inst; // @[cpu.scala 76:29]
  wire [63:0] memory_io_ex2mem_pc; // @[cpu.scala 76:29]
  wire [63:0] memory_io_ex2mem_excep_cause; // @[cpu.scala 76:29]
  wire [63:0] memory_io_ex2mem_excep_tval; // @[cpu.scala 76:29]
  wire  memory_io_ex2mem_excep_en; // @[cpu.scala 76:29]
  wire [63:0] memory_io_ex2mem_excep_pc; // @[cpu.scala 76:29]
  wire [1:0] memory_io_ex2mem_excep_etype; // @[cpu.scala 76:29]
  wire [4:0] memory_io_ex2mem_ctrl_dcMode; // @[cpu.scala 76:29]
  wire  memory_io_ex2mem_ctrl_writeRegEn; // @[cpu.scala 76:29]
  wire  memory_io_ex2mem_ctrl_writeCSREn; // @[cpu.scala 76:29]
  wire [63:0] memory_io_ex2mem_mem_addr; // @[cpu.scala 76:29]
  wire [63:0] memory_io_ex2mem_mem_data; // @[cpu.scala 76:29]
  wire [11:0] memory_io_ex2mem_csr_id; // @[cpu.scala 76:29]
  wire [63:0] memory_io_ex2mem_csr_d; // @[cpu.scala 76:29]
  wire [4:0] memory_io_ex2mem_dst; // @[cpu.scala 76:29]
  wire [63:0] memory_io_ex2mem_dst_d; // @[cpu.scala 76:29]
  wire [11:0] memory_io_ex2mem_rcsr_id; // @[cpu.scala 76:29]
  wire [1:0] memory_io_ex2mem_special; // @[cpu.scala 76:29]
  wire [1:0] memory_io_ex2mem_indi; // @[cpu.scala 76:29]
  wire  memory_io_ex2mem_drop; // @[cpu.scala 76:29]
  wire  memory_io_ex2mem_stall; // @[cpu.scala 76:29]
  wire  memory_io_ex2mem_recov; // @[cpu.scala 76:29]
  wire  memory_io_ex2mem_valid; // @[cpu.scala 76:29]
  wire  memory_io_ex2mem_ready; // @[cpu.scala 76:29]
  wire [31:0] memory_io_mem2rb_inst; // @[cpu.scala 76:29]
  wire [63:0] memory_io_mem2rb_pc; // @[cpu.scala 76:29]
  wire [63:0] memory_io_mem2rb_excep_cause; // @[cpu.scala 76:29]
  wire [63:0] memory_io_mem2rb_excep_tval; // @[cpu.scala 76:29]
  wire  memory_io_mem2rb_excep_en; // @[cpu.scala 76:29]
  wire [63:0] memory_io_mem2rb_excep_pc; // @[cpu.scala 76:29]
  wire [1:0] memory_io_mem2rb_excep_etype; // @[cpu.scala 76:29]
  wire [11:0] memory_io_mem2rb_csr_id; // @[cpu.scala 76:29]
  wire [63:0] memory_io_mem2rb_csr_d; // @[cpu.scala 76:29]
  wire  memory_io_mem2rb_csr_en; // @[cpu.scala 76:29]
  wire [4:0] memory_io_mem2rb_dst; // @[cpu.scala 76:29]
  wire [63:0] memory_io_mem2rb_dst_d; // @[cpu.scala 76:29]
  wire  memory_io_mem2rb_dst_en; // @[cpu.scala 76:29]
  wire [11:0] memory_io_mem2rb_rcsr_id; // @[cpu.scala 76:29]
  wire [1:0] memory_io_mem2rb_special; // @[cpu.scala 76:29]
  wire  memory_io_mem2rb_is_mmio; // @[cpu.scala 76:29]
  wire  memory_io_mem2rb_drop; // @[cpu.scala 76:29]
  wire  memory_io_mem2rb_stall; // @[cpu.scala 76:29]
  wire  memory_io_mem2rb_recov; // @[cpu.scala 76:29]
  wire  memory_io_mem2rb_valid; // @[cpu.scala 76:29]
  wire  memory_io_mem2rb_ready; // @[cpu.scala 76:29]
  wire [31:0] memory_io_dataRW_addr; // @[cpu.scala 76:29]
  wire [63:0] memory_io_dataRW_rdata; // @[cpu.scala 76:29]
  wire  memory_io_dataRW_rvalid; // @[cpu.scala 76:29]
  wire [63:0] memory_io_dataRW_wdata; // @[cpu.scala 76:29]
  wire [4:0] memory_io_dataRW_dc_mode; // @[cpu.scala 76:29]
  wire [4:0] memory_io_dataRW_amo; // @[cpu.scala 76:29]
  wire  memory_io_dataRW_ready; // @[cpu.scala 76:29]
  wire [63:0] memory_io_va2pa_vaddr; // @[cpu.scala 76:29]
  wire  memory_io_va2pa_vvalid; // @[cpu.scala 76:29]
  wire [1:0] memory_io_va2pa_m_type; // @[cpu.scala 76:29]
  wire [31:0] memory_io_va2pa_paddr; // @[cpu.scala 76:29]
  wire  memory_io_va2pa_pvalid; // @[cpu.scala 76:29]
  wire [63:0] memory_io_va2pa_tlb_excep_cause; // @[cpu.scala 76:29]
  wire [63:0] memory_io_va2pa_tlb_excep_tval; // @[cpu.scala 76:29]
  wire  memory_io_va2pa_tlb_excep_en; // @[cpu.scala 76:29]
  wire [4:0] memory_io_d_mem1_id; // @[cpu.scala 76:29]
  wire [63:0] memory_io_d_mem1_data; // @[cpu.scala 76:29]
  wire [1:0] memory_io_d_mem1_state; // @[cpu.scala 76:29]
  wire [4:0] memory_io_d_mem2_id; // @[cpu.scala 76:29]
  wire [63:0] memory_io_d_mem2_data; // @[cpu.scala 76:29]
  wire [1:0] memory_io_d_mem2_state; // @[cpu.scala 76:29]
  wire [4:0] memory_io_d_mem3_id; // @[cpu.scala 76:29]
  wire [63:0] memory_io_d_mem3_data; // @[cpu.scala 76:29]
  wire [1:0] memory_io_d_mem3_state; // @[cpu.scala 76:29]
  wire  writeback_clock; // @[cpu.scala 77:29]
  wire  writeback_reset; // @[cpu.scala 77:29]
  wire [31:0] writeback_io_mem2rb_inst; // @[cpu.scala 77:29]
  wire [63:0] writeback_io_mem2rb_pc; // @[cpu.scala 77:29]
  wire [63:0] writeback_io_mem2rb_excep_cause; // @[cpu.scala 77:29]
  wire [63:0] writeback_io_mem2rb_excep_tval; // @[cpu.scala 77:29]
  wire  writeback_io_mem2rb_excep_en; // @[cpu.scala 77:29]
  wire [63:0] writeback_io_mem2rb_excep_pc; // @[cpu.scala 77:29]
  wire [1:0] writeback_io_mem2rb_excep_etype; // @[cpu.scala 77:29]
  wire [11:0] writeback_io_mem2rb_csr_id; // @[cpu.scala 77:29]
  wire [63:0] writeback_io_mem2rb_csr_d; // @[cpu.scala 77:29]
  wire  writeback_io_mem2rb_csr_en; // @[cpu.scala 77:29]
  wire [4:0] writeback_io_mem2rb_dst; // @[cpu.scala 77:29]
  wire [63:0] writeback_io_mem2rb_dst_d; // @[cpu.scala 77:29]
  wire  writeback_io_mem2rb_dst_en; // @[cpu.scala 77:29]
  wire [11:0] writeback_io_mem2rb_rcsr_id; // @[cpu.scala 77:29]
  wire [1:0] writeback_io_mem2rb_special; // @[cpu.scala 77:29]
  wire  writeback_io_mem2rb_is_mmio; // @[cpu.scala 77:29]
  wire  writeback_io_mem2rb_drop; // @[cpu.scala 77:29]
  wire  writeback_io_mem2rb_stall; // @[cpu.scala 77:29]
  wire  writeback_io_mem2rb_recov; // @[cpu.scala 77:29]
  wire  writeback_io_mem2rb_valid; // @[cpu.scala 77:29]
  wire  writeback_io_mem2rb_ready; // @[cpu.scala 77:29]
  wire [4:0] writeback_io_wReg_id; // @[cpu.scala 77:29]
  wire [63:0] writeback_io_wReg_data; // @[cpu.scala 77:29]
  wire  writeback_io_wReg_en; // @[cpu.scala 77:29]
  wire [11:0] writeback_io_wCsr_id; // @[cpu.scala 77:29]
  wire [63:0] writeback_io_wCsr_data; // @[cpu.scala 77:29]
  wire  writeback_io_wCsr_en; // @[cpu.scala 77:29]
  wire [63:0] writeback_io_excep_cause; // @[cpu.scala 77:29]
  wire [63:0] writeback_io_excep_tval; // @[cpu.scala 77:29]
  wire  writeback_io_excep_en; // @[cpu.scala 77:29]
  wire [63:0] writeback_io_excep_pc; // @[cpu.scala 77:29]
  wire [1:0] writeback_io_excep_etype; // @[cpu.scala 77:29]
  wire [63:0] writeback_io_wb2if_seq_pc; // @[cpu.scala 77:29]
  wire  writeback_io_wb2if_valid; // @[cpu.scala 77:29]
  wire  writeback_io_recov; // @[cpu.scala 77:29]
  wire  writeback_io_flush_tlb; // @[cpu.scala 77:29]
  wire  writeback_io_flush_cache; // @[cpu.scala 77:29]
  wire  regs_clock; // @[cpu.scala 79:29]
  wire  regs_reset; // @[cpu.scala 79:29]
  wire [4:0] regs_io_rs1_id; // @[cpu.scala 79:29]
  wire [63:0] regs_io_rs1_data; // @[cpu.scala 79:29]
  wire [4:0] regs_io_rs2_id; // @[cpu.scala 79:29]
  wire [63:0] regs_io_rs2_data; // @[cpu.scala 79:29]
  wire [4:0] regs_io_dst_id; // @[cpu.scala 79:29]
  wire [63:0] regs_io_dst_data; // @[cpu.scala 79:29]
  wire  regs_io_dst_en; // @[cpu.scala 79:29]
  wire  csrs_clock; // @[cpu.scala 80:29]
  wire  csrs_reset; // @[cpu.scala 80:29]
  wire [11:0] csrs_io_rs_id; // @[cpu.scala 80:29]
  wire [63:0] csrs_io_rs_data; // @[cpu.scala 80:29]
  wire  csrs_io_rs_is_err; // @[cpu.scala 80:29]
  wire [11:0] csrs_io_rd_id; // @[cpu.scala 80:29]
  wire [63:0] csrs_io_rd_data; // @[cpu.scala 80:29]
  wire  csrs_io_rd_en; // @[cpu.scala 80:29]
  wire [63:0] csrs_io_excep_cause; // @[cpu.scala 80:29]
  wire [63:0] csrs_io_excep_tval; // @[cpu.scala 80:29]
  wire  csrs_io_excep_en; // @[cpu.scala 80:29]
  wire [63:0] csrs_io_excep_pc; // @[cpu.scala 80:29]
  wire [1:0] csrs_io_excep_etype; // @[cpu.scala 80:29]
  wire [1:0] csrs_io_mmuState_priv; // @[cpu.scala 80:29]
  wire [63:0] csrs_io_mmuState_mstatus; // @[cpu.scala 80:29]
  wire [63:0] csrs_io_mmuState_satp; // @[cpu.scala 80:29]
  wire [1:0] csrs_io_idState_priv; // @[cpu.scala 80:29]
  wire [63:0] csrs_io_reg2if_seq_pc; // @[cpu.scala 80:29]
  wire  csrs_io_reg2if_valid; // @[cpu.scala 80:29]
  wire  csrs_io_intr_out_en; // @[cpu.scala 80:29]
  wire [63:0] csrs_io_intr_out_cause; // @[cpu.scala 80:29]
  wire  csrs_io_clint_raise; // @[cpu.scala 80:29]
  wire  csrs_io_clint_clear; // @[cpu.scala 80:29]
  wire  csrs_io_plic_m_raise; // @[cpu.scala 80:29]
  wire  csrs_io_plic_m_clear; // @[cpu.scala 80:29]
  wire  csrs_io_plic_s_raise; // @[cpu.scala 80:29]
  wire  csrs_io_plic_s_clear; // @[cpu.scala 80:29]
  wire [63:0] csrs_io_updateNextPc_seq_pc; // @[cpu.scala 80:29]
  wire  csrs_io_updateNextPc_valid; // @[cpu.scala 80:29]
  wire  csrs_io_intr_msip_raise; // @[cpu.scala 80:29]
  wire  csrs_io_intr_msip_clear; // @[cpu.scala 80:29]
  wire  icache_clock; // @[cpu.scala 81:29]
  wire  icache_reset; // @[cpu.scala 81:29]
  wire  icache_io_instAxi_ra_ready; // @[cpu.scala 81:29]
  wire  icache_io_instAxi_ra_valid; // @[cpu.scala 81:29]
  wire [31:0] icache_io_instAxi_ra_bits_addr; // @[cpu.scala 81:29]
  wire  icache_io_instAxi_rd_valid; // @[cpu.scala 81:29]
  wire [63:0] icache_io_instAxi_rd_bits_data; // @[cpu.scala 81:29]
  wire  icache_io_instAxi_rd_bits_last; // @[cpu.scala 81:29]
  wire [31:0] icache_io_icRead_addr; // @[cpu.scala 81:29]
  wire [63:0] icache_io_icRead_inst; // @[cpu.scala 81:29]
  wire  icache_io_icRead_arvalid; // @[cpu.scala 81:29]
  wire  icache_io_icRead_ready; // @[cpu.scala 81:29]
  wire  icache_io_icRead_rvalid; // @[cpu.scala 81:29]
  wire  icache_io_flush; // @[cpu.scala 81:29]
  wire [5:0] icache_io_ic2sr0_addr; // @[cpu.scala 81:29]
  wire  icache_io_ic2sr0_cen; // @[cpu.scala 81:29]
  wire  icache_io_ic2sr0_wen; // @[cpu.scala 81:29]
  wire [127:0] icache_io_ic2sr0_wmask; // @[cpu.scala 81:29]
  wire [127:0] icache_io_ic2sr0_wdata; // @[cpu.scala 81:29]
  wire [127:0] icache_io_ic2sr0_rdata; // @[cpu.scala 81:29]
  wire [5:0] icache_io_ic2sr1_addr; // @[cpu.scala 81:29]
  wire  icache_io_ic2sr1_cen; // @[cpu.scala 81:29]
  wire  icache_io_ic2sr1_wen; // @[cpu.scala 81:29]
  wire [127:0] icache_io_ic2sr1_wmask; // @[cpu.scala 81:29]
  wire [127:0] icache_io_ic2sr1_wdata; // @[cpu.scala 81:29]
  wire [127:0] icache_io_ic2sr1_rdata; // @[cpu.scala 81:29]
  wire [5:0] icache_io_ic2sr2_addr; // @[cpu.scala 81:29]
  wire  icache_io_ic2sr2_cen; // @[cpu.scala 81:29]
  wire  icache_io_ic2sr2_wen; // @[cpu.scala 81:29]
  wire [127:0] icache_io_ic2sr2_wmask; // @[cpu.scala 81:29]
  wire [127:0] icache_io_ic2sr2_wdata; // @[cpu.scala 81:29]
  wire [127:0] icache_io_ic2sr2_rdata; // @[cpu.scala 81:29]
  wire [5:0] icache_io_ic2sr3_addr; // @[cpu.scala 81:29]
  wire  icache_io_ic2sr3_cen; // @[cpu.scala 81:29]
  wire  icache_io_ic2sr3_wen; // @[cpu.scala 81:29]
  wire [127:0] icache_io_ic2sr3_wmask; // @[cpu.scala 81:29]
  wire [127:0] icache_io_ic2sr3_wdata; // @[cpu.scala 81:29]
  wire [127:0] icache_io_ic2sr3_rdata; // @[cpu.scala 81:29]
  wire  dcache_clock; // @[cpu.scala 82:29]
  wire  dcache_reset; // @[cpu.scala 82:29]
  wire  dcache_io_dataAxi_wa_ready; // @[cpu.scala 82:29]
  wire  dcache_io_dataAxi_wa_valid; // @[cpu.scala 82:29]
  wire [31:0] dcache_io_dataAxi_wa_bits_addr; // @[cpu.scala 82:29]
  wire  dcache_io_dataAxi_wd_ready; // @[cpu.scala 82:29]
  wire  dcache_io_dataAxi_wd_valid; // @[cpu.scala 82:29]
  wire [63:0] dcache_io_dataAxi_wd_bits_data; // @[cpu.scala 82:29]
  wire  dcache_io_dataAxi_wd_bits_last; // @[cpu.scala 82:29]
  wire  dcache_io_dataAxi_ra_ready; // @[cpu.scala 82:29]
  wire  dcache_io_dataAxi_ra_valid; // @[cpu.scala 82:29]
  wire [31:0] dcache_io_dataAxi_ra_bits_addr; // @[cpu.scala 82:29]
  wire  dcache_io_dataAxi_rd_valid; // @[cpu.scala 82:29]
  wire [63:0] dcache_io_dataAxi_rd_bits_data; // @[cpu.scala 82:29]
  wire  dcache_io_dataAxi_rd_bits_last; // @[cpu.scala 82:29]
  wire [31:0] dcache_io_dcRW_addr; // @[cpu.scala 82:29]
  wire [63:0] dcache_io_dcRW_rdata; // @[cpu.scala 82:29]
  wire  dcache_io_dcRW_rvalid; // @[cpu.scala 82:29]
  wire [63:0] dcache_io_dcRW_wdata; // @[cpu.scala 82:29]
  wire [4:0] dcache_io_dcRW_dc_mode; // @[cpu.scala 82:29]
  wire [4:0] dcache_io_dcRW_amo; // @[cpu.scala 82:29]
  wire  dcache_io_dcRW_ready; // @[cpu.scala 82:29]
  wire  dcache_io_flush; // @[cpu.scala 82:29]
  wire  dcache_io_flush_out; // @[cpu.scala 82:29]
  wire [5:0] dcache_io_dc2sr0_addr; // @[cpu.scala 82:29]
  wire  dcache_io_dc2sr0_cen; // @[cpu.scala 82:29]
  wire  dcache_io_dc2sr0_wen; // @[cpu.scala 82:29]
  wire [127:0] dcache_io_dc2sr0_wmask; // @[cpu.scala 82:29]
  wire [127:0] dcache_io_dc2sr0_wdata; // @[cpu.scala 82:29]
  wire [127:0] dcache_io_dc2sr0_rdata; // @[cpu.scala 82:29]
  wire [5:0] dcache_io_dc2sr1_addr; // @[cpu.scala 82:29]
  wire  dcache_io_dc2sr1_cen; // @[cpu.scala 82:29]
  wire  dcache_io_dc2sr1_wen; // @[cpu.scala 82:29]
  wire [127:0] dcache_io_dc2sr1_wmask; // @[cpu.scala 82:29]
  wire [127:0] dcache_io_dc2sr1_wdata; // @[cpu.scala 82:29]
  wire [127:0] dcache_io_dc2sr1_rdata; // @[cpu.scala 82:29]
  wire [5:0] dcache_io_dc2sr2_addr; // @[cpu.scala 82:29]
  wire  dcache_io_dc2sr2_cen; // @[cpu.scala 82:29]
  wire  dcache_io_dc2sr2_wen; // @[cpu.scala 82:29]
  wire [127:0] dcache_io_dc2sr2_wmask; // @[cpu.scala 82:29]
  wire [127:0] dcache_io_dc2sr2_wdata; // @[cpu.scala 82:29]
  wire [127:0] dcache_io_dc2sr2_rdata; // @[cpu.scala 82:29]
  wire [5:0] dcache_io_dc2sr3_addr; // @[cpu.scala 82:29]
  wire  dcache_io_dc2sr3_cen; // @[cpu.scala 82:29]
  wire  dcache_io_dc2sr3_wen; // @[cpu.scala 82:29]
  wire [127:0] dcache_io_dc2sr3_wmask; // @[cpu.scala 82:29]
  wire [127:0] dcache_io_dc2sr3_wdata; // @[cpu.scala 82:29]
  wire [127:0] dcache_io_dc2sr3_rdata; // @[cpu.scala 82:29]
  wire  mem2Axi_clock; // @[cpu.scala 84:29]
  wire  mem2Axi_reset; // @[cpu.scala 84:29]
  wire [31:0] mem2Axi_io_dataIO_addr; // @[cpu.scala 84:29]
  wire [63:0] mem2Axi_io_dataIO_rdata; // @[cpu.scala 84:29]
  wire  mem2Axi_io_dataIO_rvalid; // @[cpu.scala 84:29]
  wire [63:0] mem2Axi_io_dataIO_wdata; // @[cpu.scala 84:29]
  wire [4:0] mem2Axi_io_dataIO_dc_mode; // @[cpu.scala 84:29]
  wire  mem2Axi_io_dataIO_ready; // @[cpu.scala 84:29]
  wire  mem2Axi_io_outAxi_wa_ready; // @[cpu.scala 84:29]
  wire  mem2Axi_io_outAxi_wa_valid; // @[cpu.scala 84:29]
  wire [3:0] mem2Axi_io_outAxi_wa_bits_id; // @[cpu.scala 84:29]
  wire [31:0] mem2Axi_io_outAxi_wa_bits_addr; // @[cpu.scala 84:29]
  wire [7:0] mem2Axi_io_outAxi_wa_bits_len; // @[cpu.scala 84:29]
  wire [2:0] mem2Axi_io_outAxi_wa_bits_size; // @[cpu.scala 84:29]
  wire [1:0] mem2Axi_io_outAxi_wa_bits_burst; // @[cpu.scala 84:29]
  wire  mem2Axi_io_outAxi_wd_ready; // @[cpu.scala 84:29]
  wire  mem2Axi_io_outAxi_wd_valid; // @[cpu.scala 84:29]
  wire [63:0] mem2Axi_io_outAxi_wd_bits_data; // @[cpu.scala 84:29]
  wire [7:0] mem2Axi_io_outAxi_wd_bits_strb; // @[cpu.scala 84:29]
  wire  mem2Axi_io_outAxi_wd_bits_last; // @[cpu.scala 84:29]
  wire  mem2Axi_io_outAxi_wr_ready; // @[cpu.scala 84:29]
  wire  mem2Axi_io_outAxi_wr_valid; // @[cpu.scala 84:29]
  wire [3:0] mem2Axi_io_outAxi_wr_bits_id; // @[cpu.scala 84:29]
  wire [1:0] mem2Axi_io_outAxi_wr_bits_resp; // @[cpu.scala 84:29]
  wire  mem2Axi_io_outAxi_ra_ready; // @[cpu.scala 84:29]
  wire  mem2Axi_io_outAxi_ra_valid; // @[cpu.scala 84:29]
  wire [3:0] mem2Axi_io_outAxi_ra_bits_id; // @[cpu.scala 84:29]
  wire [31:0] mem2Axi_io_outAxi_ra_bits_addr; // @[cpu.scala 84:29]
  wire [7:0] mem2Axi_io_outAxi_ra_bits_len; // @[cpu.scala 84:29]
  wire [2:0] mem2Axi_io_outAxi_ra_bits_size; // @[cpu.scala 84:29]
  wire [1:0] mem2Axi_io_outAxi_ra_bits_burst; // @[cpu.scala 84:29]
  wire  mem2Axi_io_outAxi_rd_ready; // @[cpu.scala 84:29]
  wire  mem2Axi_io_outAxi_rd_valid; // @[cpu.scala 84:29]
  wire [3:0] mem2Axi_io_outAxi_rd_bits_id; // @[cpu.scala 84:29]
  wire [63:0] mem2Axi_io_outAxi_rd_bits_data; // @[cpu.scala 84:29]
  wire [1:0] mem2Axi_io_outAxi_rd_bits_resp; // @[cpu.scala 84:29]
  wire  mem2Axi_io_outAxi_rd_bits_last; // @[cpu.scala 84:29]
  wire  flash2Axi_clock; // @[cpu.scala 85:29]
  wire  flash2Axi_reset; // @[cpu.scala 85:29]
  wire [31:0] flash2Axi_io_dataIO_addr; // @[cpu.scala 85:29]
  wire [63:0] flash2Axi_io_dataIO_rdata; // @[cpu.scala 85:29]
  wire  flash2Axi_io_dataIO_rvalid; // @[cpu.scala 85:29]
  wire [63:0] flash2Axi_io_dataIO_wdata; // @[cpu.scala 85:29]
  wire [4:0] flash2Axi_io_dataIO_dc_mode; // @[cpu.scala 85:29]
  wire  flash2Axi_io_dataIO_ready; // @[cpu.scala 85:29]
  wire  flash2Axi_io_outAxi_wa_ready; // @[cpu.scala 85:29]
  wire  flash2Axi_io_outAxi_wa_valid; // @[cpu.scala 85:29]
  wire [3:0] flash2Axi_io_outAxi_wa_bits_id; // @[cpu.scala 85:29]
  wire [31:0] flash2Axi_io_outAxi_wa_bits_addr; // @[cpu.scala 85:29]
  wire [7:0] flash2Axi_io_outAxi_wa_bits_len; // @[cpu.scala 85:29]
  wire [2:0] flash2Axi_io_outAxi_wa_bits_size; // @[cpu.scala 85:29]
  wire [1:0] flash2Axi_io_outAxi_wa_bits_burst; // @[cpu.scala 85:29]
  wire  flash2Axi_io_outAxi_wd_ready; // @[cpu.scala 85:29]
  wire  flash2Axi_io_outAxi_wd_valid; // @[cpu.scala 85:29]
  wire [63:0] flash2Axi_io_outAxi_wd_bits_data; // @[cpu.scala 85:29]
  wire [7:0] flash2Axi_io_outAxi_wd_bits_strb; // @[cpu.scala 85:29]
  wire  flash2Axi_io_outAxi_wd_bits_last; // @[cpu.scala 85:29]
  wire  flash2Axi_io_outAxi_wr_ready; // @[cpu.scala 85:29]
  wire  flash2Axi_io_outAxi_wr_valid; // @[cpu.scala 85:29]
  wire [3:0] flash2Axi_io_outAxi_wr_bits_id; // @[cpu.scala 85:29]
  wire [1:0] flash2Axi_io_outAxi_wr_bits_resp; // @[cpu.scala 85:29]
  wire  flash2Axi_io_outAxi_ra_ready; // @[cpu.scala 85:29]
  wire  flash2Axi_io_outAxi_ra_valid; // @[cpu.scala 85:29]
  wire [3:0] flash2Axi_io_outAxi_ra_bits_id; // @[cpu.scala 85:29]
  wire [31:0] flash2Axi_io_outAxi_ra_bits_addr; // @[cpu.scala 85:29]
  wire [7:0] flash2Axi_io_outAxi_ra_bits_len; // @[cpu.scala 85:29]
  wire [2:0] flash2Axi_io_outAxi_ra_bits_size; // @[cpu.scala 85:29]
  wire [1:0] flash2Axi_io_outAxi_ra_bits_burst; // @[cpu.scala 85:29]
  wire  flash2Axi_io_outAxi_rd_ready; // @[cpu.scala 85:29]
  wire  flash2Axi_io_outAxi_rd_valid; // @[cpu.scala 85:29]
  wire [3:0] flash2Axi_io_outAxi_rd_bits_id; // @[cpu.scala 85:29]
  wire [63:0] flash2Axi_io_outAxi_rd_bits_data; // @[cpu.scala 85:29]
  wire [1:0] flash2Axi_io_outAxi_rd_bits_resp; // @[cpu.scala 85:29]
  wire  flash2Axi_io_outAxi_rd_bits_last; // @[cpu.scala 85:29]
  wire  crossBar_clock; // @[cpu.scala 87:29]
  wire  crossBar_reset; // @[cpu.scala 87:29]
  wire  crossBar_io_icAxi_ra_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_icAxi_ra_valid; // @[cpu.scala 87:29]
  wire [31:0] crossBar_io_icAxi_ra_bits_addr; // @[cpu.scala 87:29]
  wire  crossBar_io_icAxi_rd_valid; // @[cpu.scala 87:29]
  wire [63:0] crossBar_io_icAxi_rd_bits_data; // @[cpu.scala 87:29]
  wire  crossBar_io_icAxi_rd_bits_last; // @[cpu.scala 87:29]
  wire  crossBar_io_flashAxi_wa_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_flashAxi_wa_valid; // @[cpu.scala 87:29]
  wire [3:0] crossBar_io_flashAxi_wa_bits_id; // @[cpu.scala 87:29]
  wire [31:0] crossBar_io_flashAxi_wa_bits_addr; // @[cpu.scala 87:29]
  wire [7:0] crossBar_io_flashAxi_wa_bits_len; // @[cpu.scala 87:29]
  wire [2:0] crossBar_io_flashAxi_wa_bits_size; // @[cpu.scala 87:29]
  wire [1:0] crossBar_io_flashAxi_wa_bits_burst; // @[cpu.scala 87:29]
  wire  crossBar_io_flashAxi_wd_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_flashAxi_wd_valid; // @[cpu.scala 87:29]
  wire [63:0] crossBar_io_flashAxi_wd_bits_data; // @[cpu.scala 87:29]
  wire [7:0] crossBar_io_flashAxi_wd_bits_strb; // @[cpu.scala 87:29]
  wire  crossBar_io_flashAxi_wd_bits_last; // @[cpu.scala 87:29]
  wire  crossBar_io_flashAxi_wr_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_flashAxi_wr_valid; // @[cpu.scala 87:29]
  wire [3:0] crossBar_io_flashAxi_wr_bits_id; // @[cpu.scala 87:29]
  wire [1:0] crossBar_io_flashAxi_wr_bits_resp; // @[cpu.scala 87:29]
  wire  crossBar_io_flashAxi_ra_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_flashAxi_ra_valid; // @[cpu.scala 87:29]
  wire [3:0] crossBar_io_flashAxi_ra_bits_id; // @[cpu.scala 87:29]
  wire [31:0] crossBar_io_flashAxi_ra_bits_addr; // @[cpu.scala 87:29]
  wire [7:0] crossBar_io_flashAxi_ra_bits_len; // @[cpu.scala 87:29]
  wire [2:0] crossBar_io_flashAxi_ra_bits_size; // @[cpu.scala 87:29]
  wire [1:0] crossBar_io_flashAxi_ra_bits_burst; // @[cpu.scala 87:29]
  wire  crossBar_io_flashAxi_rd_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_flashAxi_rd_valid; // @[cpu.scala 87:29]
  wire [3:0] crossBar_io_flashAxi_rd_bits_id; // @[cpu.scala 87:29]
  wire [63:0] crossBar_io_flashAxi_rd_bits_data; // @[cpu.scala 87:29]
  wire [1:0] crossBar_io_flashAxi_rd_bits_resp; // @[cpu.scala 87:29]
  wire  crossBar_io_flashAxi_rd_bits_last; // @[cpu.scala 87:29]
  wire  crossBar_io_memAxi_wa_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_memAxi_wa_valid; // @[cpu.scala 87:29]
  wire [31:0] crossBar_io_memAxi_wa_bits_addr; // @[cpu.scala 87:29]
  wire  crossBar_io_memAxi_wd_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_memAxi_wd_valid; // @[cpu.scala 87:29]
  wire [63:0] crossBar_io_memAxi_wd_bits_data; // @[cpu.scala 87:29]
  wire  crossBar_io_memAxi_wd_bits_last; // @[cpu.scala 87:29]
  wire  crossBar_io_memAxi_ra_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_memAxi_ra_valid; // @[cpu.scala 87:29]
  wire [31:0] crossBar_io_memAxi_ra_bits_addr; // @[cpu.scala 87:29]
  wire  crossBar_io_memAxi_rd_valid; // @[cpu.scala 87:29]
  wire [63:0] crossBar_io_memAxi_rd_bits_data; // @[cpu.scala 87:29]
  wire  crossBar_io_memAxi_rd_bits_last; // @[cpu.scala 87:29]
  wire  crossBar_io_mmioAxi_wa_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_mmioAxi_wa_valid; // @[cpu.scala 87:29]
  wire [3:0] crossBar_io_mmioAxi_wa_bits_id; // @[cpu.scala 87:29]
  wire [31:0] crossBar_io_mmioAxi_wa_bits_addr; // @[cpu.scala 87:29]
  wire [7:0] crossBar_io_mmioAxi_wa_bits_len; // @[cpu.scala 87:29]
  wire [2:0] crossBar_io_mmioAxi_wa_bits_size; // @[cpu.scala 87:29]
  wire [1:0] crossBar_io_mmioAxi_wa_bits_burst; // @[cpu.scala 87:29]
  wire  crossBar_io_mmioAxi_wd_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_mmioAxi_wd_valid; // @[cpu.scala 87:29]
  wire [63:0] crossBar_io_mmioAxi_wd_bits_data; // @[cpu.scala 87:29]
  wire [7:0] crossBar_io_mmioAxi_wd_bits_strb; // @[cpu.scala 87:29]
  wire  crossBar_io_mmioAxi_wd_bits_last; // @[cpu.scala 87:29]
  wire  crossBar_io_mmioAxi_wr_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_mmioAxi_wr_valid; // @[cpu.scala 87:29]
  wire [3:0] crossBar_io_mmioAxi_wr_bits_id; // @[cpu.scala 87:29]
  wire [1:0] crossBar_io_mmioAxi_wr_bits_resp; // @[cpu.scala 87:29]
  wire  crossBar_io_mmioAxi_ra_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_mmioAxi_ra_valid; // @[cpu.scala 87:29]
  wire [3:0] crossBar_io_mmioAxi_ra_bits_id; // @[cpu.scala 87:29]
  wire [31:0] crossBar_io_mmioAxi_ra_bits_addr; // @[cpu.scala 87:29]
  wire [7:0] crossBar_io_mmioAxi_ra_bits_len; // @[cpu.scala 87:29]
  wire [2:0] crossBar_io_mmioAxi_ra_bits_size; // @[cpu.scala 87:29]
  wire [1:0] crossBar_io_mmioAxi_ra_bits_burst; // @[cpu.scala 87:29]
  wire  crossBar_io_mmioAxi_rd_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_mmioAxi_rd_valid; // @[cpu.scala 87:29]
  wire [3:0] crossBar_io_mmioAxi_rd_bits_id; // @[cpu.scala 87:29]
  wire [63:0] crossBar_io_mmioAxi_rd_bits_data; // @[cpu.scala 87:29]
  wire [1:0] crossBar_io_mmioAxi_rd_bits_resp; // @[cpu.scala 87:29]
  wire  crossBar_io_mmioAxi_rd_bits_last; // @[cpu.scala 87:29]
  wire  crossBar_io_outAxi_wa_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_outAxi_wa_valid; // @[cpu.scala 87:29]
  wire [3:0] crossBar_io_outAxi_wa_bits_id; // @[cpu.scala 87:29]
  wire [31:0] crossBar_io_outAxi_wa_bits_addr; // @[cpu.scala 87:29]
  wire [7:0] crossBar_io_outAxi_wa_bits_len; // @[cpu.scala 87:29]
  wire [2:0] crossBar_io_outAxi_wa_bits_size; // @[cpu.scala 87:29]
  wire [1:0] crossBar_io_outAxi_wa_bits_burst; // @[cpu.scala 87:29]
  wire  crossBar_io_outAxi_wd_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_outAxi_wd_valid; // @[cpu.scala 87:29]
  wire [63:0] crossBar_io_outAxi_wd_bits_data; // @[cpu.scala 87:29]
  wire [7:0] crossBar_io_outAxi_wd_bits_strb; // @[cpu.scala 87:29]
  wire  crossBar_io_outAxi_wd_bits_last; // @[cpu.scala 87:29]
  wire  crossBar_io_outAxi_wr_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_outAxi_wr_valid; // @[cpu.scala 87:29]
  wire [3:0] crossBar_io_outAxi_wr_bits_id; // @[cpu.scala 87:29]
  wire [1:0] crossBar_io_outAxi_wr_bits_resp; // @[cpu.scala 87:29]
  wire  crossBar_io_outAxi_ra_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_outAxi_ra_valid; // @[cpu.scala 87:29]
  wire [3:0] crossBar_io_outAxi_ra_bits_id; // @[cpu.scala 87:29]
  wire [31:0] crossBar_io_outAxi_ra_bits_addr; // @[cpu.scala 87:29]
  wire [7:0] crossBar_io_outAxi_ra_bits_len; // @[cpu.scala 87:29]
  wire [2:0] crossBar_io_outAxi_ra_bits_size; // @[cpu.scala 87:29]
  wire [1:0] crossBar_io_outAxi_ra_bits_burst; // @[cpu.scala 87:29]
  wire  crossBar_io_outAxi_rd_ready; // @[cpu.scala 87:29]
  wire  crossBar_io_outAxi_rd_valid; // @[cpu.scala 87:29]
  wire [3:0] crossBar_io_outAxi_rd_bits_id; // @[cpu.scala 87:29]
  wire [63:0] crossBar_io_outAxi_rd_bits_data; // @[cpu.scala 87:29]
  wire [1:0] crossBar_io_outAxi_rd_bits_resp; // @[cpu.scala 87:29]
  wire  crossBar_io_outAxi_rd_bits_last; // @[cpu.scala 87:29]
  wire  crossBar_io_selectMem; // @[cpu.scala 87:29]
  wire  fetchCrossbar_clock; // @[cpu.scala 88:31]
  wire  fetchCrossbar_reset; // @[cpu.scala 88:31]
  wire [31:0] fetchCrossbar_io_instIO_addr; // @[cpu.scala 88:31]
  wire [63:0] fetchCrossbar_io_instIO_inst; // @[cpu.scala 88:31]
  wire  fetchCrossbar_io_instIO_arvalid; // @[cpu.scala 88:31]
  wire  fetchCrossbar_io_instIO_rvalid; // @[cpu.scala 88:31]
  wire [31:0] fetchCrossbar_io_icRead_addr; // @[cpu.scala 88:31]
  wire [63:0] fetchCrossbar_io_icRead_inst; // @[cpu.scala 88:31]
  wire  fetchCrossbar_io_icRead_arvalid; // @[cpu.scala 88:31]
  wire  fetchCrossbar_io_icRead_rvalid; // @[cpu.scala 88:31]
  wire [31:0] fetchCrossbar_io_flashRead_addr; // @[cpu.scala 88:31]
  wire [63:0] fetchCrossbar_io_flashRead_rdata; // @[cpu.scala 88:31]
  wire  fetchCrossbar_io_flashRead_rvalid; // @[cpu.scala 88:31]
  wire [4:0] fetchCrossbar_io_flashRead_dc_mode; // @[cpu.scala 88:31]
  wire  split64to32_clock; // @[cpu.scala 89:29]
  wire  split64to32_reset; // @[cpu.scala 89:29]
  wire [31:0] split64to32_io_data_in_addr; // @[cpu.scala 89:29]
  wire [63:0] split64to32_io_data_in_rdata; // @[cpu.scala 89:29]
  wire  split64to32_io_data_in_rvalid; // @[cpu.scala 89:29]
  wire [4:0] split64to32_io_data_in_dc_mode; // @[cpu.scala 89:29]
  wire [31:0] split64to32_io_data_out_addr; // @[cpu.scala 89:29]
  wire [63:0] split64to32_io_data_out_rdata; // @[cpu.scala 89:29]
  wire  split64to32_io_data_out_rvalid; // @[cpu.scala 89:29]
  wire [4:0] split64to32_io_data_out_dc_mode; // @[cpu.scala 89:29]
  wire  split64to32_io_data_out_ready; // @[cpu.scala 89:29]
  wire  memCrossbar_clock; // @[cpu.scala 90:29]
  wire  memCrossbar_reset; // @[cpu.scala 90:29]
  wire [31:0] memCrossbar_io_dataRW_addr; // @[cpu.scala 90:29]
  wire [63:0] memCrossbar_io_dataRW_rdata; // @[cpu.scala 90:29]
  wire  memCrossbar_io_dataRW_rvalid; // @[cpu.scala 90:29]
  wire [63:0] memCrossbar_io_dataRW_wdata; // @[cpu.scala 90:29]
  wire [4:0] memCrossbar_io_dataRW_dc_mode; // @[cpu.scala 90:29]
  wire [4:0] memCrossbar_io_dataRW_amo; // @[cpu.scala 90:29]
  wire  memCrossbar_io_dataRW_ready; // @[cpu.scala 90:29]
  wire [31:0] memCrossbar_io_mmio_addr; // @[cpu.scala 90:29]
  wire [63:0] memCrossbar_io_mmio_rdata; // @[cpu.scala 90:29]
  wire  memCrossbar_io_mmio_rvalid; // @[cpu.scala 90:29]
  wire [63:0] memCrossbar_io_mmio_wdata; // @[cpu.scala 90:29]
  wire [4:0] memCrossbar_io_mmio_dc_mode; // @[cpu.scala 90:29]
  wire  memCrossbar_io_mmio_ready; // @[cpu.scala 90:29]
  wire [31:0] memCrossbar_io_dcRW_addr; // @[cpu.scala 90:29]
  wire [63:0] memCrossbar_io_dcRW_rdata; // @[cpu.scala 90:29]
  wire  memCrossbar_io_dcRW_rvalid; // @[cpu.scala 90:29]
  wire [63:0] memCrossbar_io_dcRW_wdata; // @[cpu.scala 90:29]
  wire [4:0] memCrossbar_io_dcRW_dc_mode; // @[cpu.scala 90:29]
  wire [4:0] memCrossbar_io_dcRW_amo; // @[cpu.scala 90:29]
  wire  memCrossbar_io_dcRW_ready; // @[cpu.scala 90:29]
  wire [31:0] memCrossbar_io_clintIO_addr; // @[cpu.scala 90:29]
  wire [63:0] memCrossbar_io_clintIO_rdata; // @[cpu.scala 90:29]
  wire [63:0] memCrossbar_io_clintIO_wdata; // @[cpu.scala 90:29]
  wire  memCrossbar_io_clintIO_wvalid; // @[cpu.scala 90:29]
  wire [31:0] memCrossbar_io_plicIO_addr; // @[cpu.scala 90:29]
  wire [63:0] memCrossbar_io_plicIO_rdata; // @[cpu.scala 90:29]
  wire [63:0] memCrossbar_io_plicIO_wdata; // @[cpu.scala 90:29]
  wire  memCrossbar_io_plicIO_wvalid; // @[cpu.scala 90:29]
  wire  memCrossbar_io_plicIO_arvalid; // @[cpu.scala 90:29]
  wire  tlb_if_clock; // @[cpu.scala 91:30]
  wire  tlb_if_reset; // @[cpu.scala 91:30]
  wire [63:0] tlb_if_io_va2pa_vaddr; // @[cpu.scala 91:30]
  wire  tlb_if_io_va2pa_vvalid; // @[cpu.scala 91:30]
  wire  tlb_if_io_va2pa_ready; // @[cpu.scala 91:30]
  wire [31:0] tlb_if_io_va2pa_paddr; // @[cpu.scala 91:30]
  wire  tlb_if_io_va2pa_pvalid; // @[cpu.scala 91:30]
  wire [63:0] tlb_if_io_va2pa_tlb_excep_cause; // @[cpu.scala 91:30]
  wire [63:0] tlb_if_io_va2pa_tlb_excep_tval; // @[cpu.scala 91:30]
  wire  tlb_if_io_va2pa_tlb_excep_en; // @[cpu.scala 91:30]
  wire [1:0] tlb_if_io_mmuState_priv; // @[cpu.scala 91:30]
  wire [63:0] tlb_if_io_mmuState_mstatus; // @[cpu.scala 91:30]
  wire [63:0] tlb_if_io_mmuState_satp; // @[cpu.scala 91:30]
  wire  tlb_if_io_flush; // @[cpu.scala 91:30]
  wire [31:0] tlb_if_io_dcacheRW_addr; // @[cpu.scala 91:30]
  wire [63:0] tlb_if_io_dcacheRW_rdata; // @[cpu.scala 91:30]
  wire  tlb_if_io_dcacheRW_rvalid; // @[cpu.scala 91:30]
  wire [63:0] tlb_if_io_dcacheRW_wdata; // @[cpu.scala 91:30]
  wire [4:0] tlb_if_io_dcacheRW_dc_mode; // @[cpu.scala 91:30]
  wire  tlb_if_io_dcacheRW_ready; // @[cpu.scala 91:30]
  wire  tlb_mem_clock; // @[cpu.scala 92:30]
  wire  tlb_mem_reset; // @[cpu.scala 92:30]
  wire [63:0] tlb_mem_io_va2pa_vaddr; // @[cpu.scala 92:30]
  wire  tlb_mem_io_va2pa_vvalid; // @[cpu.scala 92:30]
  wire [1:0] tlb_mem_io_va2pa_m_type; // @[cpu.scala 92:30]
  wire  tlb_mem_io_va2pa_ready; // @[cpu.scala 92:30]
  wire [31:0] tlb_mem_io_va2pa_paddr; // @[cpu.scala 92:30]
  wire  tlb_mem_io_va2pa_pvalid; // @[cpu.scala 92:30]
  wire [63:0] tlb_mem_io_va2pa_tlb_excep_cause; // @[cpu.scala 92:30]
  wire [63:0] tlb_mem_io_va2pa_tlb_excep_tval; // @[cpu.scala 92:30]
  wire  tlb_mem_io_va2pa_tlb_excep_en; // @[cpu.scala 92:30]
  wire [1:0] tlb_mem_io_mmuState_priv; // @[cpu.scala 92:30]
  wire [63:0] tlb_mem_io_mmuState_mstatus; // @[cpu.scala 92:30]
  wire [63:0] tlb_mem_io_mmuState_satp; // @[cpu.scala 92:30]
  wire  tlb_mem_io_flush; // @[cpu.scala 92:30]
  wire [31:0] tlb_mem_io_dcacheRW_addr; // @[cpu.scala 92:30]
  wire [63:0] tlb_mem_io_dcacheRW_rdata; // @[cpu.scala 92:30]
  wire  tlb_mem_io_dcacheRW_rvalid; // @[cpu.scala 92:30]
  wire [63:0] tlb_mem_io_dcacheRW_wdata; // @[cpu.scala 92:30]
  wire [4:0] tlb_mem_io_dcacheRW_dc_mode; // @[cpu.scala 92:30]
  wire  tlb_mem_io_dcacheRW_ready; // @[cpu.scala 92:30]
  wire  dcSelector_clock; // @[cpu.scala 93:29]
  wire  dcSelector_reset; // @[cpu.scala 93:29]
  wire [31:0] dcSelector_io_tlb_if2dc_addr; // @[cpu.scala 93:29]
  wire [63:0] dcSelector_io_tlb_if2dc_rdata; // @[cpu.scala 93:29]
  wire  dcSelector_io_tlb_if2dc_rvalid; // @[cpu.scala 93:29]
  wire [63:0] dcSelector_io_tlb_if2dc_wdata; // @[cpu.scala 93:29]
  wire [4:0] dcSelector_io_tlb_if2dc_dc_mode; // @[cpu.scala 93:29]
  wire  dcSelector_io_tlb_if2dc_ready; // @[cpu.scala 93:29]
  wire [31:0] dcSelector_io_tlb_mem2dc_addr; // @[cpu.scala 93:29]
  wire [63:0] dcSelector_io_tlb_mem2dc_rdata; // @[cpu.scala 93:29]
  wire  dcSelector_io_tlb_mem2dc_rvalid; // @[cpu.scala 93:29]
  wire [63:0] dcSelector_io_tlb_mem2dc_wdata; // @[cpu.scala 93:29]
  wire [4:0] dcSelector_io_tlb_mem2dc_dc_mode; // @[cpu.scala 93:29]
  wire  dcSelector_io_tlb_mem2dc_ready; // @[cpu.scala 93:29]
  wire [31:0] dcSelector_io_mem2dc_addr; // @[cpu.scala 93:29]
  wire [63:0] dcSelector_io_mem2dc_rdata; // @[cpu.scala 93:29]
  wire  dcSelector_io_mem2dc_rvalid; // @[cpu.scala 93:29]
  wire [63:0] dcSelector_io_mem2dc_wdata; // @[cpu.scala 93:29]
  wire [4:0] dcSelector_io_mem2dc_dc_mode; // @[cpu.scala 93:29]
  wire [4:0] dcSelector_io_mem2dc_amo; // @[cpu.scala 93:29]
  wire  dcSelector_io_mem2dc_ready; // @[cpu.scala 93:29]
  wire [31:0] dcSelector_io_dma2dc_addr; // @[cpu.scala 93:29]
  wire [63:0] dcSelector_io_dma2dc_rdata; // @[cpu.scala 93:29]
  wire  dcSelector_io_dma2dc_rvalid; // @[cpu.scala 93:29]
  wire [63:0] dcSelector_io_dma2dc_wdata; // @[cpu.scala 93:29]
  wire [4:0] dcSelector_io_dma2dc_dc_mode; // @[cpu.scala 93:29]
  wire  dcSelector_io_dma2dc_ready; // @[cpu.scala 93:29]
  wire [31:0] dcSelector_io_select_addr; // @[cpu.scala 93:29]
  wire [63:0] dcSelector_io_select_rdata; // @[cpu.scala 93:29]
  wire  dcSelector_io_select_rvalid; // @[cpu.scala 93:29]
  wire [63:0] dcSelector_io_select_wdata; // @[cpu.scala 93:29]
  wire [4:0] dcSelector_io_select_dc_mode; // @[cpu.scala 93:29]
  wire [4:0] dcSelector_io_select_amo; // @[cpu.scala 93:29]
  wire  dcSelector_io_select_ready; // @[cpu.scala 93:29]
  wire  clint_clock; // @[cpu.scala 94:29]
  wire  clint_reset; // @[cpu.scala 94:29]
  wire [31:0] clint_io_rw_addr; // @[cpu.scala 94:29]
  wire [63:0] clint_io_rw_rdata; // @[cpu.scala 94:29]
  wire [63:0] clint_io_rw_wdata; // @[cpu.scala 94:29]
  wire  clint_io_rw_wvalid; // @[cpu.scala 94:29]
  wire  clint_io_intr_raise; // @[cpu.scala 94:29]
  wire  clint_io_intr_clear; // @[cpu.scala 94:29]
  wire  clint_io_intr_msip_raise; // @[cpu.scala 94:29]
  wire  clint_io_intr_msip_clear; // @[cpu.scala 94:29]
  wire  plic_clock; // @[cpu.scala 95:29]
  wire  plic_reset; // @[cpu.scala 95:29]
  wire  plic_io_intr_in1; // @[cpu.scala 95:29]
  wire  plic_io_intr_out_m_raise; // @[cpu.scala 95:29]
  wire  plic_io_intr_out_m_clear; // @[cpu.scala 95:29]
  wire  plic_io_intr_out_s_raise; // @[cpu.scala 95:29]
  wire  plic_io_intr_out_s_clear; // @[cpu.scala 95:29]
  wire [31:0] plic_io_rw_addr; // @[cpu.scala 95:29]
  wire [63:0] plic_io_rw_rdata; // @[cpu.scala 95:29]
  wire [63:0] plic_io_rw_wdata; // @[cpu.scala 95:29]
  wire  plic_io_rw_wvalid; // @[cpu.scala 95:29]
  wire  plic_io_rw_arvalid; // @[cpu.scala 95:29]
  wire  dmaBridge_clock; // @[cpu.scala 96:29]
  wire  dmaBridge_reset; // @[cpu.scala 96:29]
  wire  dmaBridge_io_dmaAxi_awready; // @[cpu.scala 96:29]
  wire  dmaBridge_io_dmaAxi_awvalid; // @[cpu.scala 96:29]
  wire [31:0] dmaBridge_io_dmaAxi_awaddr; // @[cpu.scala 96:29]
  wire [3:0] dmaBridge_io_dmaAxi_awid; // @[cpu.scala 96:29]
  wire [7:0] dmaBridge_io_dmaAxi_awlen; // @[cpu.scala 96:29]
  wire [2:0] dmaBridge_io_dmaAxi_awsize; // @[cpu.scala 96:29]
  wire  dmaBridge_io_dmaAxi_wready; // @[cpu.scala 96:29]
  wire  dmaBridge_io_dmaAxi_wvalid; // @[cpu.scala 96:29]
  wire [63:0] dmaBridge_io_dmaAxi_wdata; // @[cpu.scala 96:29]
  wire [7:0] dmaBridge_io_dmaAxi_wstrb; // @[cpu.scala 96:29]
  wire  dmaBridge_io_dmaAxi_bready; // @[cpu.scala 96:29]
  wire  dmaBridge_io_dmaAxi_bvalid; // @[cpu.scala 96:29]
  wire [3:0] dmaBridge_io_dmaAxi_bid; // @[cpu.scala 96:29]
  wire  dmaBridge_io_dmaAxi_arready; // @[cpu.scala 96:29]
  wire  dmaBridge_io_dmaAxi_arvalid; // @[cpu.scala 96:29]
  wire [31:0] dmaBridge_io_dmaAxi_araddr; // @[cpu.scala 96:29]
  wire [3:0] dmaBridge_io_dmaAxi_arid; // @[cpu.scala 96:29]
  wire [7:0] dmaBridge_io_dmaAxi_arlen; // @[cpu.scala 96:29]
  wire [2:0] dmaBridge_io_dmaAxi_arsize; // @[cpu.scala 96:29]
  wire  dmaBridge_io_dmaAxi_rready; // @[cpu.scala 96:29]
  wire  dmaBridge_io_dmaAxi_rvalid; // @[cpu.scala 96:29]
  wire [63:0] dmaBridge_io_dmaAxi_rdata; // @[cpu.scala 96:29]
  wire  dmaBridge_io_dmaAxi_rlast; // @[cpu.scala 96:29]
  wire [3:0] dmaBridge_io_dmaAxi_rid; // @[cpu.scala 96:29]
  wire [31:0] dmaBridge_io_dcRW_addr; // @[cpu.scala 96:29]
  wire [63:0] dmaBridge_io_dcRW_rdata; // @[cpu.scala 96:29]
  wire  dmaBridge_io_dcRW_rvalid; // @[cpu.scala 96:29]
  wire [63:0] dmaBridge_io_dcRW_wdata; // @[cpu.scala 96:29]
  wire [4:0] dmaBridge_io_dcRW_dc_mode; // @[cpu.scala 96:29]
  wire  dmaBridge_io_dcRW_ready; // @[cpu.scala 96:29]
  ysyx_210539_Fetch fetch ( // @[cpu.scala 71:29]
    .clock(fetch_clock),
    .reset(fetch_reset),
    .io_instRead_addr(fetch_io_instRead_addr),
    .io_instRead_inst(fetch_io_instRead_inst),
    .io_instRead_arvalid(fetch_io_instRead_arvalid),
    .io_instRead_rvalid(fetch_io_instRead_rvalid),
    .io_va2pa_vaddr(fetch_io_va2pa_vaddr),
    .io_va2pa_vvalid(fetch_io_va2pa_vvalid),
    .io_va2pa_paddr(fetch_io_va2pa_paddr),
    .io_va2pa_pvalid(fetch_io_va2pa_pvalid),
    .io_va2pa_tlb_excep_cause(fetch_io_va2pa_tlb_excep_cause),
    .io_va2pa_tlb_excep_tval(fetch_io_va2pa_tlb_excep_tval),
    .io_va2pa_tlb_excep_en(fetch_io_va2pa_tlb_excep_en),
    .io_reg2if_seq_pc(fetch_io_reg2if_seq_pc),
    .io_reg2if_valid(fetch_io_reg2if_valid),
    .io_wb2if_seq_pc(fetch_io_wb2if_seq_pc),
    .io_wb2if_valid(fetch_io_wb2if_valid),
    .io_recov(fetch_io_recov),
    .io_intr_in_en(fetch_io_intr_in_en),
    .io_intr_in_cause(fetch_io_intr_in_cause),
    .io_branchFail_seq_pc(fetch_io_branchFail_seq_pc),
    .io_branchFail_valid(fetch_io_branchFail_valid),
    .io_if2id_inst(fetch_io_if2id_inst),
    .io_if2id_pc(fetch_io_if2id_pc),
    .io_if2id_excep_cause(fetch_io_if2id_excep_cause),
    .io_if2id_excep_tval(fetch_io_if2id_excep_tval),
    .io_if2id_excep_en(fetch_io_if2id_excep_en),
    .io_if2id_excep_pc(fetch_io_if2id_excep_pc),
    .io_if2id_drop(fetch_io_if2id_drop),
    .io_if2id_stall(fetch_io_if2id_stall),
    .io_if2id_recov(fetch_io_if2id_recov),
    .io_if2id_valid(fetch_io_if2id_valid),
    .io_if2id_ready(fetch_io_if2id_ready)
  );
  ysyx_210539_Decode decode ( // @[cpu.scala 72:29]
    .clock(decode_clock),
    .reset(decode_reset),
    .io_if2id_inst(decode_io_if2id_inst),
    .io_if2id_pc(decode_io_if2id_pc),
    .io_if2id_excep_cause(decode_io_if2id_excep_cause),
    .io_if2id_excep_tval(decode_io_if2id_excep_tval),
    .io_if2id_excep_en(decode_io_if2id_excep_en),
    .io_if2id_excep_pc(decode_io_if2id_excep_pc),
    .io_if2id_drop(decode_io_if2id_drop),
    .io_if2id_stall(decode_io_if2id_stall),
    .io_if2id_recov(decode_io_if2id_recov),
    .io_if2id_valid(decode_io_if2id_valid),
    .io_if2id_ready(decode_io_if2id_ready),
    .io_id2df_inst(decode_io_id2df_inst),
    .io_id2df_pc(decode_io_id2df_pc),
    .io_id2df_excep_cause(decode_io_id2df_excep_cause),
    .io_id2df_excep_tval(decode_io_id2df_excep_tval),
    .io_id2df_excep_en(decode_io_id2df_excep_en),
    .io_id2df_excep_pc(decode_io_id2df_excep_pc),
    .io_id2df_excep_etype(decode_io_id2df_excep_etype),
    .io_id2df_ctrl_aluOp(decode_io_id2df_ctrl_aluOp),
    .io_id2df_ctrl_aluWidth(decode_io_id2df_ctrl_aluWidth),
    .io_id2df_ctrl_dcMode(decode_io_id2df_ctrl_dcMode),
    .io_id2df_ctrl_writeRegEn(decode_io_id2df_ctrl_writeRegEn),
    .io_id2df_ctrl_writeCSREn(decode_io_id2df_ctrl_writeCSREn),
    .io_id2df_ctrl_brType(decode_io_id2df_ctrl_brType),
    .io_id2df_rs1(decode_io_id2df_rs1),
    .io_id2df_rrs1(decode_io_id2df_rrs1),
    .io_id2df_rs1_d(decode_io_id2df_rs1_d),
    .io_id2df_rs2(decode_io_id2df_rs2),
    .io_id2df_rrs2(decode_io_id2df_rrs2),
    .io_id2df_rs2_d(decode_io_id2df_rs2_d),
    .io_id2df_dst(decode_io_id2df_dst),
    .io_id2df_dst_d(decode_io_id2df_dst_d),
    .io_id2df_jmp_type(decode_io_id2df_jmp_type),
    .io_id2df_special(decode_io_id2df_special),
    .io_id2df_swap(decode_io_id2df_swap),
    .io_id2df_indi(decode_io_id2df_indi),
    .io_id2df_drop(decode_io_id2df_drop),
    .io_id2df_stall(decode_io_id2df_stall),
    .io_id2df_recov(decode_io_id2df_recov),
    .io_id2df_valid(decode_io_id2df_valid),
    .io_id2df_ready(decode_io_id2df_ready),
    .io_idState_priv(decode_io_idState_priv)
  );
  ysyx_210539_Forwarding forwading ( // @[cpu.scala 73:29]
    .clock(forwading_clock),
    .reset(forwading_reset),
    .io_id2df_inst(forwading_io_id2df_inst),
    .io_id2df_pc(forwading_io_id2df_pc),
    .io_id2df_excep_cause(forwading_io_id2df_excep_cause),
    .io_id2df_excep_tval(forwading_io_id2df_excep_tval),
    .io_id2df_excep_en(forwading_io_id2df_excep_en),
    .io_id2df_excep_pc(forwading_io_id2df_excep_pc),
    .io_id2df_excep_etype(forwading_io_id2df_excep_etype),
    .io_id2df_ctrl_aluOp(forwading_io_id2df_ctrl_aluOp),
    .io_id2df_ctrl_aluWidth(forwading_io_id2df_ctrl_aluWidth),
    .io_id2df_ctrl_dcMode(forwading_io_id2df_ctrl_dcMode),
    .io_id2df_ctrl_writeRegEn(forwading_io_id2df_ctrl_writeRegEn),
    .io_id2df_ctrl_writeCSREn(forwading_io_id2df_ctrl_writeCSREn),
    .io_id2df_ctrl_brType(forwading_io_id2df_ctrl_brType),
    .io_id2df_rs1(forwading_io_id2df_rs1),
    .io_id2df_rrs1(forwading_io_id2df_rrs1),
    .io_id2df_rs1_d(forwading_io_id2df_rs1_d),
    .io_id2df_rs2(forwading_io_id2df_rs2),
    .io_id2df_rrs2(forwading_io_id2df_rrs2),
    .io_id2df_rs2_d(forwading_io_id2df_rs2_d),
    .io_id2df_dst(forwading_io_id2df_dst),
    .io_id2df_dst_d(forwading_io_id2df_dst_d),
    .io_id2df_jmp_type(forwading_io_id2df_jmp_type),
    .io_id2df_special(forwading_io_id2df_special),
    .io_id2df_swap(forwading_io_id2df_swap),
    .io_id2df_indi(forwading_io_id2df_indi),
    .io_id2df_drop(forwading_io_id2df_drop),
    .io_id2df_stall(forwading_io_id2df_stall),
    .io_id2df_recov(forwading_io_id2df_recov),
    .io_id2df_valid(forwading_io_id2df_valid),
    .io_id2df_ready(forwading_io_id2df_ready),
    .io_df2rr_inst(forwading_io_df2rr_inst),
    .io_df2rr_pc(forwading_io_df2rr_pc),
    .io_df2rr_excep_cause(forwading_io_df2rr_excep_cause),
    .io_df2rr_excep_tval(forwading_io_df2rr_excep_tval),
    .io_df2rr_excep_en(forwading_io_df2rr_excep_en),
    .io_df2rr_excep_pc(forwading_io_df2rr_excep_pc),
    .io_df2rr_excep_etype(forwading_io_df2rr_excep_etype),
    .io_df2rr_ctrl_aluOp(forwading_io_df2rr_ctrl_aluOp),
    .io_df2rr_ctrl_aluWidth(forwading_io_df2rr_ctrl_aluWidth),
    .io_df2rr_ctrl_dcMode(forwading_io_df2rr_ctrl_dcMode),
    .io_df2rr_ctrl_writeRegEn(forwading_io_df2rr_ctrl_writeRegEn),
    .io_df2rr_ctrl_writeCSREn(forwading_io_df2rr_ctrl_writeCSREn),
    .io_df2rr_ctrl_brType(forwading_io_df2rr_ctrl_brType),
    .io_df2rr_rs1(forwading_io_df2rr_rs1),
    .io_df2rr_rrs1(forwading_io_df2rr_rrs1),
    .io_df2rr_rs1_d(forwading_io_df2rr_rs1_d),
    .io_df2rr_rs2(forwading_io_df2rr_rs2),
    .io_df2rr_rrs2(forwading_io_df2rr_rrs2),
    .io_df2rr_rs2_d(forwading_io_df2rr_rs2_d),
    .io_df2rr_dst(forwading_io_df2rr_dst),
    .io_df2rr_dst_d(forwading_io_df2rr_dst_d),
    .io_df2rr_jmp_type(forwading_io_df2rr_jmp_type),
    .io_df2rr_special(forwading_io_df2rr_special),
    .io_df2rr_swap(forwading_io_df2rr_swap),
    .io_df2rr_indi(forwading_io_df2rr_indi),
    .io_df2rr_drop(forwading_io_df2rr_drop),
    .io_df2rr_stall(forwading_io_df2rr_stall),
    .io_df2rr_recov(forwading_io_df2rr_recov),
    .io_df2rr_valid(forwading_io_df2rr_valid),
    .io_df2rr_ready(forwading_io_df2rr_ready),
    .io_d_rr_id(forwading_io_d_rr_id),
    .io_d_rr_data(forwading_io_d_rr_data),
    .io_d_rr_state(forwading_io_d_rr_state),
    .io_d_ex_id(forwading_io_d_ex_id),
    .io_d_ex_data(forwading_io_d_ex_data),
    .io_d_ex_state(forwading_io_d_ex_state),
    .io_d_mem1_id(forwading_io_d_mem1_id),
    .io_d_mem1_data(forwading_io_d_mem1_data),
    .io_d_mem1_state(forwading_io_d_mem1_state),
    .io_d_mem2_id(forwading_io_d_mem2_id),
    .io_d_mem2_data(forwading_io_d_mem2_data),
    .io_d_mem2_state(forwading_io_d_mem2_state),
    .io_d_mem3_id(forwading_io_d_mem3_id),
    .io_d_mem3_data(forwading_io_d_mem3_data),
    .io_d_mem3_state(forwading_io_d_mem3_state)
  );
  ysyx_210539_ReadRegs readregs ( // @[cpu.scala 74:29]
    .clock(readregs_clock),
    .reset(readregs_reset),
    .io_df2rr_inst(readregs_io_df2rr_inst),
    .io_df2rr_pc(readregs_io_df2rr_pc),
    .io_df2rr_excep_cause(readregs_io_df2rr_excep_cause),
    .io_df2rr_excep_tval(readregs_io_df2rr_excep_tval),
    .io_df2rr_excep_en(readregs_io_df2rr_excep_en),
    .io_df2rr_excep_pc(readregs_io_df2rr_excep_pc),
    .io_df2rr_excep_etype(readregs_io_df2rr_excep_etype),
    .io_df2rr_ctrl_aluOp(readregs_io_df2rr_ctrl_aluOp),
    .io_df2rr_ctrl_aluWidth(readregs_io_df2rr_ctrl_aluWidth),
    .io_df2rr_ctrl_dcMode(readregs_io_df2rr_ctrl_dcMode),
    .io_df2rr_ctrl_writeRegEn(readregs_io_df2rr_ctrl_writeRegEn),
    .io_df2rr_ctrl_writeCSREn(readregs_io_df2rr_ctrl_writeCSREn),
    .io_df2rr_ctrl_brType(readregs_io_df2rr_ctrl_brType),
    .io_df2rr_rs1(readregs_io_df2rr_rs1),
    .io_df2rr_rrs1(readregs_io_df2rr_rrs1),
    .io_df2rr_rs1_d(readregs_io_df2rr_rs1_d),
    .io_df2rr_rs2(readregs_io_df2rr_rs2),
    .io_df2rr_rrs2(readregs_io_df2rr_rrs2),
    .io_df2rr_rs2_d(readregs_io_df2rr_rs2_d),
    .io_df2rr_dst(readregs_io_df2rr_dst),
    .io_df2rr_dst_d(readregs_io_df2rr_dst_d),
    .io_df2rr_jmp_type(readregs_io_df2rr_jmp_type),
    .io_df2rr_special(readregs_io_df2rr_special),
    .io_df2rr_swap(readregs_io_df2rr_swap),
    .io_df2rr_indi(readregs_io_df2rr_indi),
    .io_df2rr_drop(readregs_io_df2rr_drop),
    .io_df2rr_stall(readregs_io_df2rr_stall),
    .io_df2rr_recov(readregs_io_df2rr_recov),
    .io_df2rr_valid(readregs_io_df2rr_valid),
    .io_df2rr_ready(readregs_io_df2rr_ready),
    .io_rr2ex_inst(readregs_io_rr2ex_inst),
    .io_rr2ex_pc(readregs_io_rr2ex_pc),
    .io_rr2ex_excep_cause(readregs_io_rr2ex_excep_cause),
    .io_rr2ex_excep_tval(readregs_io_rr2ex_excep_tval),
    .io_rr2ex_excep_en(readregs_io_rr2ex_excep_en),
    .io_rr2ex_excep_pc(readregs_io_rr2ex_excep_pc),
    .io_rr2ex_excep_etype(readregs_io_rr2ex_excep_etype),
    .io_rr2ex_ctrl_aluOp(readregs_io_rr2ex_ctrl_aluOp),
    .io_rr2ex_ctrl_aluWidth(readregs_io_rr2ex_ctrl_aluWidth),
    .io_rr2ex_ctrl_dcMode(readregs_io_rr2ex_ctrl_dcMode),
    .io_rr2ex_ctrl_writeRegEn(readregs_io_rr2ex_ctrl_writeRegEn),
    .io_rr2ex_ctrl_writeCSREn(readregs_io_rr2ex_ctrl_writeCSREn),
    .io_rr2ex_ctrl_brType(readregs_io_rr2ex_ctrl_brType),
    .io_rr2ex_rs1_d(readregs_io_rr2ex_rs1_d),
    .io_rr2ex_rs2(readregs_io_rr2ex_rs2),
    .io_rr2ex_rs2_d(readregs_io_rr2ex_rs2_d),
    .io_rr2ex_dst(readregs_io_rr2ex_dst),
    .io_rr2ex_dst_d(readregs_io_rr2ex_dst_d),
    .io_rr2ex_rcsr_id(readregs_io_rr2ex_rcsr_id),
    .io_rr2ex_jmp_type(readregs_io_rr2ex_jmp_type),
    .io_rr2ex_special(readregs_io_rr2ex_special),
    .io_rr2ex_indi(readregs_io_rr2ex_indi),
    .io_rr2ex_drop(readregs_io_rr2ex_drop),
    .io_rr2ex_stall(readregs_io_rr2ex_stall),
    .io_rr2ex_recov(readregs_io_rr2ex_recov),
    .io_rr2ex_valid(readregs_io_rr2ex_valid),
    .io_rr2ex_ready(readregs_io_rr2ex_ready),
    .io_rs1Read_id(readregs_io_rs1Read_id),
    .io_rs1Read_data(readregs_io_rs1Read_data),
    .io_rs2Read_id(readregs_io_rs2Read_id),
    .io_rs2Read_data(readregs_io_rs2Read_data),
    .io_csrRead_id(readregs_io_csrRead_id),
    .io_csrRead_data(readregs_io_csrRead_data),
    .io_csrRead_is_err(readregs_io_csrRead_is_err),
    .io_d_rr_id(readregs_io_d_rr_id),
    .io_d_rr_data(readregs_io_d_rr_data),
    .io_d_rr_state(readregs_io_d_rr_state)
  );
  ysyx_210539_Execute execute ( // @[cpu.scala 75:29]
    .clock(execute_clock),
    .reset(execute_reset),
    .io_rr2ex_inst(execute_io_rr2ex_inst),
    .io_rr2ex_pc(execute_io_rr2ex_pc),
    .io_rr2ex_excep_cause(execute_io_rr2ex_excep_cause),
    .io_rr2ex_excep_tval(execute_io_rr2ex_excep_tval),
    .io_rr2ex_excep_en(execute_io_rr2ex_excep_en),
    .io_rr2ex_excep_pc(execute_io_rr2ex_excep_pc),
    .io_rr2ex_excep_etype(execute_io_rr2ex_excep_etype),
    .io_rr2ex_ctrl_aluOp(execute_io_rr2ex_ctrl_aluOp),
    .io_rr2ex_ctrl_aluWidth(execute_io_rr2ex_ctrl_aluWidth),
    .io_rr2ex_ctrl_dcMode(execute_io_rr2ex_ctrl_dcMode),
    .io_rr2ex_ctrl_writeRegEn(execute_io_rr2ex_ctrl_writeRegEn),
    .io_rr2ex_ctrl_writeCSREn(execute_io_rr2ex_ctrl_writeCSREn),
    .io_rr2ex_ctrl_brType(execute_io_rr2ex_ctrl_brType),
    .io_rr2ex_rs1_d(execute_io_rr2ex_rs1_d),
    .io_rr2ex_rs2(execute_io_rr2ex_rs2),
    .io_rr2ex_rs2_d(execute_io_rr2ex_rs2_d),
    .io_rr2ex_dst(execute_io_rr2ex_dst),
    .io_rr2ex_dst_d(execute_io_rr2ex_dst_d),
    .io_rr2ex_rcsr_id(execute_io_rr2ex_rcsr_id),
    .io_rr2ex_jmp_type(execute_io_rr2ex_jmp_type),
    .io_rr2ex_special(execute_io_rr2ex_special),
    .io_rr2ex_indi(execute_io_rr2ex_indi),
    .io_rr2ex_drop(execute_io_rr2ex_drop),
    .io_rr2ex_stall(execute_io_rr2ex_stall),
    .io_rr2ex_recov(execute_io_rr2ex_recov),
    .io_rr2ex_valid(execute_io_rr2ex_valid),
    .io_rr2ex_ready(execute_io_rr2ex_ready),
    .io_ex2mem_inst(execute_io_ex2mem_inst),
    .io_ex2mem_pc(execute_io_ex2mem_pc),
    .io_ex2mem_excep_cause(execute_io_ex2mem_excep_cause),
    .io_ex2mem_excep_tval(execute_io_ex2mem_excep_tval),
    .io_ex2mem_excep_en(execute_io_ex2mem_excep_en),
    .io_ex2mem_excep_pc(execute_io_ex2mem_excep_pc),
    .io_ex2mem_excep_etype(execute_io_ex2mem_excep_etype),
    .io_ex2mem_ctrl_dcMode(execute_io_ex2mem_ctrl_dcMode),
    .io_ex2mem_ctrl_writeRegEn(execute_io_ex2mem_ctrl_writeRegEn),
    .io_ex2mem_ctrl_writeCSREn(execute_io_ex2mem_ctrl_writeCSREn),
    .io_ex2mem_mem_addr(execute_io_ex2mem_mem_addr),
    .io_ex2mem_mem_data(execute_io_ex2mem_mem_data),
    .io_ex2mem_csr_id(execute_io_ex2mem_csr_id),
    .io_ex2mem_csr_d(execute_io_ex2mem_csr_d),
    .io_ex2mem_dst(execute_io_ex2mem_dst),
    .io_ex2mem_dst_d(execute_io_ex2mem_dst_d),
    .io_ex2mem_rcsr_id(execute_io_ex2mem_rcsr_id),
    .io_ex2mem_special(execute_io_ex2mem_special),
    .io_ex2mem_indi(execute_io_ex2mem_indi),
    .io_ex2mem_drop(execute_io_ex2mem_drop),
    .io_ex2mem_stall(execute_io_ex2mem_stall),
    .io_ex2mem_recov(execute_io_ex2mem_recov),
    .io_ex2mem_valid(execute_io_ex2mem_valid),
    .io_ex2mem_ready(execute_io_ex2mem_ready),
    .io_d_ex_id(execute_io_d_ex_id),
    .io_d_ex_data(execute_io_d_ex_data),
    .io_d_ex_state(execute_io_d_ex_state),
    .io_ex2if_seq_pc(execute_io_ex2if_seq_pc),
    .io_ex2if_valid(execute_io_ex2if_valid),
    .io_updateNextPc_seq_pc(execute_io_updateNextPc_seq_pc),
    .io_updateNextPc_valid(execute_io_updateNextPc_valid)
  );
  ysyx_210539_Memory memory ( // @[cpu.scala 76:29]
    .clock(memory_clock),
    .reset(memory_reset),
    .io_ex2mem_inst(memory_io_ex2mem_inst),
    .io_ex2mem_pc(memory_io_ex2mem_pc),
    .io_ex2mem_excep_cause(memory_io_ex2mem_excep_cause),
    .io_ex2mem_excep_tval(memory_io_ex2mem_excep_tval),
    .io_ex2mem_excep_en(memory_io_ex2mem_excep_en),
    .io_ex2mem_excep_pc(memory_io_ex2mem_excep_pc),
    .io_ex2mem_excep_etype(memory_io_ex2mem_excep_etype),
    .io_ex2mem_ctrl_dcMode(memory_io_ex2mem_ctrl_dcMode),
    .io_ex2mem_ctrl_writeRegEn(memory_io_ex2mem_ctrl_writeRegEn),
    .io_ex2mem_ctrl_writeCSREn(memory_io_ex2mem_ctrl_writeCSREn),
    .io_ex2mem_mem_addr(memory_io_ex2mem_mem_addr),
    .io_ex2mem_mem_data(memory_io_ex2mem_mem_data),
    .io_ex2mem_csr_id(memory_io_ex2mem_csr_id),
    .io_ex2mem_csr_d(memory_io_ex2mem_csr_d),
    .io_ex2mem_dst(memory_io_ex2mem_dst),
    .io_ex2mem_dst_d(memory_io_ex2mem_dst_d),
    .io_ex2mem_rcsr_id(memory_io_ex2mem_rcsr_id),
    .io_ex2mem_special(memory_io_ex2mem_special),
    .io_ex2mem_indi(memory_io_ex2mem_indi),
    .io_ex2mem_drop(memory_io_ex2mem_drop),
    .io_ex2mem_stall(memory_io_ex2mem_stall),
    .io_ex2mem_recov(memory_io_ex2mem_recov),
    .io_ex2mem_valid(memory_io_ex2mem_valid),
    .io_ex2mem_ready(memory_io_ex2mem_ready),
    .io_mem2rb_inst(memory_io_mem2rb_inst),
    .io_mem2rb_pc(memory_io_mem2rb_pc),
    .io_mem2rb_excep_cause(memory_io_mem2rb_excep_cause),
    .io_mem2rb_excep_tval(memory_io_mem2rb_excep_tval),
    .io_mem2rb_excep_en(memory_io_mem2rb_excep_en),
    .io_mem2rb_excep_pc(memory_io_mem2rb_excep_pc),
    .io_mem2rb_excep_etype(memory_io_mem2rb_excep_etype),
    .io_mem2rb_csr_id(memory_io_mem2rb_csr_id),
    .io_mem2rb_csr_d(memory_io_mem2rb_csr_d),
    .io_mem2rb_csr_en(memory_io_mem2rb_csr_en),
    .io_mem2rb_dst(memory_io_mem2rb_dst),
    .io_mem2rb_dst_d(memory_io_mem2rb_dst_d),
    .io_mem2rb_dst_en(memory_io_mem2rb_dst_en),
    .io_mem2rb_rcsr_id(memory_io_mem2rb_rcsr_id),
    .io_mem2rb_special(memory_io_mem2rb_special),
    .io_mem2rb_is_mmio(memory_io_mem2rb_is_mmio),
    .io_mem2rb_drop(memory_io_mem2rb_drop),
    .io_mem2rb_stall(memory_io_mem2rb_stall),
    .io_mem2rb_recov(memory_io_mem2rb_recov),
    .io_mem2rb_valid(memory_io_mem2rb_valid),
    .io_mem2rb_ready(memory_io_mem2rb_ready),
    .io_dataRW_addr(memory_io_dataRW_addr),
    .io_dataRW_rdata(memory_io_dataRW_rdata),
    .io_dataRW_rvalid(memory_io_dataRW_rvalid),
    .io_dataRW_wdata(memory_io_dataRW_wdata),
    .io_dataRW_dc_mode(memory_io_dataRW_dc_mode),
    .io_dataRW_amo(memory_io_dataRW_amo),
    .io_dataRW_ready(memory_io_dataRW_ready),
    .io_va2pa_vaddr(memory_io_va2pa_vaddr),
    .io_va2pa_vvalid(memory_io_va2pa_vvalid),
    .io_va2pa_m_type(memory_io_va2pa_m_type),
    .io_va2pa_paddr(memory_io_va2pa_paddr),
    .io_va2pa_pvalid(memory_io_va2pa_pvalid),
    .io_va2pa_tlb_excep_cause(memory_io_va2pa_tlb_excep_cause),
    .io_va2pa_tlb_excep_tval(memory_io_va2pa_tlb_excep_tval),
    .io_va2pa_tlb_excep_en(memory_io_va2pa_tlb_excep_en),
    .io_d_mem1_id(memory_io_d_mem1_id),
    .io_d_mem1_data(memory_io_d_mem1_data),
    .io_d_mem1_state(memory_io_d_mem1_state),
    .io_d_mem2_id(memory_io_d_mem2_id),
    .io_d_mem2_data(memory_io_d_mem2_data),
    .io_d_mem2_state(memory_io_d_mem2_state),
    .io_d_mem3_id(memory_io_d_mem3_id),
    .io_d_mem3_data(memory_io_d_mem3_data),
    .io_d_mem3_state(memory_io_d_mem3_state)
  );
  ysyx_210539_Writeback writeback ( // @[cpu.scala 77:29]
    .clock(writeback_clock),
    .reset(writeback_reset),
    .io_mem2rb_inst(writeback_io_mem2rb_inst),
    .io_mem2rb_pc(writeback_io_mem2rb_pc),
    .io_mem2rb_excep_cause(writeback_io_mem2rb_excep_cause),
    .io_mem2rb_excep_tval(writeback_io_mem2rb_excep_tval),
    .io_mem2rb_excep_en(writeback_io_mem2rb_excep_en),
    .io_mem2rb_excep_pc(writeback_io_mem2rb_excep_pc),
    .io_mem2rb_excep_etype(writeback_io_mem2rb_excep_etype),
    .io_mem2rb_csr_id(writeback_io_mem2rb_csr_id),
    .io_mem2rb_csr_d(writeback_io_mem2rb_csr_d),
    .io_mem2rb_csr_en(writeback_io_mem2rb_csr_en),
    .io_mem2rb_dst(writeback_io_mem2rb_dst),
    .io_mem2rb_dst_d(writeback_io_mem2rb_dst_d),
    .io_mem2rb_dst_en(writeback_io_mem2rb_dst_en),
    .io_mem2rb_rcsr_id(writeback_io_mem2rb_rcsr_id),
    .io_mem2rb_special(writeback_io_mem2rb_special),
    .io_mem2rb_is_mmio(writeback_io_mem2rb_is_mmio),
    .io_mem2rb_drop(writeback_io_mem2rb_drop),
    .io_mem2rb_stall(writeback_io_mem2rb_stall),
    .io_mem2rb_recov(writeback_io_mem2rb_recov),
    .io_mem2rb_valid(writeback_io_mem2rb_valid),
    .io_mem2rb_ready(writeback_io_mem2rb_ready),
    .io_wReg_id(writeback_io_wReg_id),
    .io_wReg_data(writeback_io_wReg_data),
    .io_wReg_en(writeback_io_wReg_en),
    .io_wCsr_id(writeback_io_wCsr_id),
    .io_wCsr_data(writeback_io_wCsr_data),
    .io_wCsr_en(writeback_io_wCsr_en),
    .io_excep_cause(writeback_io_excep_cause),
    .io_excep_tval(writeback_io_excep_tval),
    .io_excep_en(writeback_io_excep_en),
    .io_excep_pc(writeback_io_excep_pc),
    .io_excep_etype(writeback_io_excep_etype),
    .io_wb2if_seq_pc(writeback_io_wb2if_seq_pc),
    .io_wb2if_valid(writeback_io_wb2if_valid),
    .io_recov(writeback_io_recov),
    .io_flush_tlb(writeback_io_flush_tlb),
    .io_flush_cache(writeback_io_flush_cache)
  );
  ysyx_210539_Regs regs ( // @[cpu.scala 79:29]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_rs1_id(regs_io_rs1_id),
    .io_rs1_data(regs_io_rs1_data),
    .io_rs2_id(regs_io_rs2_id),
    .io_rs2_data(regs_io_rs2_data),
    .io_dst_id(regs_io_dst_id),
    .io_dst_data(regs_io_dst_data),
    .io_dst_en(regs_io_dst_en)
  );
  ysyx_210539_Csrs csrs ( // @[cpu.scala 80:29]
    .clock(csrs_clock),
    .reset(csrs_reset),
    .io_rs_id(csrs_io_rs_id),
    .io_rs_data(csrs_io_rs_data),
    .io_rs_is_err(csrs_io_rs_is_err),
    .io_rd_id(csrs_io_rd_id),
    .io_rd_data(csrs_io_rd_data),
    .io_rd_en(csrs_io_rd_en),
    .io_excep_cause(csrs_io_excep_cause),
    .io_excep_tval(csrs_io_excep_tval),
    .io_excep_en(csrs_io_excep_en),
    .io_excep_pc(csrs_io_excep_pc),
    .io_excep_etype(csrs_io_excep_etype),
    .io_mmuState_priv(csrs_io_mmuState_priv),
    .io_mmuState_mstatus(csrs_io_mmuState_mstatus),
    .io_mmuState_satp(csrs_io_mmuState_satp),
    .io_idState_priv(csrs_io_idState_priv),
    .io_reg2if_seq_pc(csrs_io_reg2if_seq_pc),
    .io_reg2if_valid(csrs_io_reg2if_valid),
    .io_intr_out_en(csrs_io_intr_out_en),
    .io_intr_out_cause(csrs_io_intr_out_cause),
    .io_clint_raise(csrs_io_clint_raise),
    .io_clint_clear(csrs_io_clint_clear),
    .io_plic_m_raise(csrs_io_plic_m_raise),
    .io_plic_m_clear(csrs_io_plic_m_clear),
    .io_plic_s_raise(csrs_io_plic_s_raise),
    .io_plic_s_clear(csrs_io_plic_s_clear),
    .io_updateNextPc_seq_pc(csrs_io_updateNextPc_seq_pc),
    .io_updateNextPc_valid(csrs_io_updateNextPc_valid),
    .io_intr_msip_raise(csrs_io_intr_msip_raise),
    .io_intr_msip_clear(csrs_io_intr_msip_clear)
  );
  ysyx_210539_InstCache icache ( // @[cpu.scala 81:29]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_instAxi_ra_ready(icache_io_instAxi_ra_ready),
    .io_instAxi_ra_valid(icache_io_instAxi_ra_valid),
    .io_instAxi_ra_bits_addr(icache_io_instAxi_ra_bits_addr),
    .io_instAxi_rd_valid(icache_io_instAxi_rd_valid),
    .io_instAxi_rd_bits_data(icache_io_instAxi_rd_bits_data),
    .io_instAxi_rd_bits_last(icache_io_instAxi_rd_bits_last),
    .io_icRead_addr(icache_io_icRead_addr),
    .io_icRead_inst(icache_io_icRead_inst),
    .io_icRead_arvalid(icache_io_icRead_arvalid),
    .io_icRead_ready(icache_io_icRead_ready),
    .io_icRead_rvalid(icache_io_icRead_rvalid),
    .io_flush(icache_io_flush),
    .io_ic2sr0_addr(icache_io_ic2sr0_addr),
    .io_ic2sr0_cen(icache_io_ic2sr0_cen),
    .io_ic2sr0_wen(icache_io_ic2sr0_wen),
    .io_ic2sr0_wmask(icache_io_ic2sr0_wmask),
    .io_ic2sr0_wdata(icache_io_ic2sr0_wdata),
    .io_ic2sr0_rdata(icache_io_ic2sr0_rdata),
    .io_ic2sr1_addr(icache_io_ic2sr1_addr),
    .io_ic2sr1_cen(icache_io_ic2sr1_cen),
    .io_ic2sr1_wen(icache_io_ic2sr1_wen),
    .io_ic2sr1_wmask(icache_io_ic2sr1_wmask),
    .io_ic2sr1_wdata(icache_io_ic2sr1_wdata),
    .io_ic2sr1_rdata(icache_io_ic2sr1_rdata),
    .io_ic2sr2_addr(icache_io_ic2sr2_addr),
    .io_ic2sr2_cen(icache_io_ic2sr2_cen),
    .io_ic2sr2_wen(icache_io_ic2sr2_wen),
    .io_ic2sr2_wmask(icache_io_ic2sr2_wmask),
    .io_ic2sr2_wdata(icache_io_ic2sr2_wdata),
    .io_ic2sr2_rdata(icache_io_ic2sr2_rdata),
    .io_ic2sr3_addr(icache_io_ic2sr3_addr),
    .io_ic2sr3_cen(icache_io_ic2sr3_cen),
    .io_ic2sr3_wen(icache_io_ic2sr3_wen),
    .io_ic2sr3_wmask(icache_io_ic2sr3_wmask),
    .io_ic2sr3_wdata(icache_io_ic2sr3_wdata),
    .io_ic2sr3_rdata(icache_io_ic2sr3_rdata)
  );
  ysyx_210539_DataCache dcache ( // @[cpu.scala 82:29]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_dataAxi_wa_ready(dcache_io_dataAxi_wa_ready),
    .io_dataAxi_wa_valid(dcache_io_dataAxi_wa_valid),
    .io_dataAxi_wa_bits_addr(dcache_io_dataAxi_wa_bits_addr),
    .io_dataAxi_wd_ready(dcache_io_dataAxi_wd_ready),
    .io_dataAxi_wd_valid(dcache_io_dataAxi_wd_valid),
    .io_dataAxi_wd_bits_data(dcache_io_dataAxi_wd_bits_data),
    .io_dataAxi_wd_bits_last(dcache_io_dataAxi_wd_bits_last),
    .io_dataAxi_ra_ready(dcache_io_dataAxi_ra_ready),
    .io_dataAxi_ra_valid(dcache_io_dataAxi_ra_valid),
    .io_dataAxi_ra_bits_addr(dcache_io_dataAxi_ra_bits_addr),
    .io_dataAxi_rd_valid(dcache_io_dataAxi_rd_valid),
    .io_dataAxi_rd_bits_data(dcache_io_dataAxi_rd_bits_data),
    .io_dataAxi_rd_bits_last(dcache_io_dataAxi_rd_bits_last),
    .io_dcRW_addr(dcache_io_dcRW_addr),
    .io_dcRW_rdata(dcache_io_dcRW_rdata),
    .io_dcRW_rvalid(dcache_io_dcRW_rvalid),
    .io_dcRW_wdata(dcache_io_dcRW_wdata),
    .io_dcRW_dc_mode(dcache_io_dcRW_dc_mode),
    .io_dcRW_amo(dcache_io_dcRW_amo),
    .io_dcRW_ready(dcache_io_dcRW_ready),
    .io_flush(dcache_io_flush),
    .io_flush_out(dcache_io_flush_out),
    .io_dc2sr0_addr(dcache_io_dc2sr0_addr),
    .io_dc2sr0_cen(dcache_io_dc2sr0_cen),
    .io_dc2sr0_wen(dcache_io_dc2sr0_wen),
    .io_dc2sr0_wmask(dcache_io_dc2sr0_wmask),
    .io_dc2sr0_wdata(dcache_io_dc2sr0_wdata),
    .io_dc2sr0_rdata(dcache_io_dc2sr0_rdata),
    .io_dc2sr1_addr(dcache_io_dc2sr1_addr),
    .io_dc2sr1_cen(dcache_io_dc2sr1_cen),
    .io_dc2sr1_wen(dcache_io_dc2sr1_wen),
    .io_dc2sr1_wmask(dcache_io_dc2sr1_wmask),
    .io_dc2sr1_wdata(dcache_io_dc2sr1_wdata),
    .io_dc2sr1_rdata(dcache_io_dc2sr1_rdata),
    .io_dc2sr2_addr(dcache_io_dc2sr2_addr),
    .io_dc2sr2_cen(dcache_io_dc2sr2_cen),
    .io_dc2sr2_wen(dcache_io_dc2sr2_wen),
    .io_dc2sr2_wmask(dcache_io_dc2sr2_wmask),
    .io_dc2sr2_wdata(dcache_io_dc2sr2_wdata),
    .io_dc2sr2_rdata(dcache_io_dc2sr2_rdata),
    .io_dc2sr3_addr(dcache_io_dc2sr3_addr),
    .io_dc2sr3_cen(dcache_io_dc2sr3_cen),
    .io_dc2sr3_wen(dcache_io_dc2sr3_wen),
    .io_dc2sr3_wmask(dcache_io_dc2sr3_wmask),
    .io_dc2sr3_wdata(dcache_io_dc2sr3_wdata),
    .io_dc2sr3_rdata(dcache_io_dc2sr3_rdata)
  );
  ysyx_210539_ToAXI mem2Axi ( // @[cpu.scala 84:29]
    .clock(mem2Axi_clock),
    .reset(mem2Axi_reset),
    .io_dataIO_addr(mem2Axi_io_dataIO_addr),
    .io_dataIO_rdata(mem2Axi_io_dataIO_rdata),
    .io_dataIO_rvalid(mem2Axi_io_dataIO_rvalid),
    .io_dataIO_wdata(mem2Axi_io_dataIO_wdata),
    .io_dataIO_dc_mode(mem2Axi_io_dataIO_dc_mode),
    .io_dataIO_ready(mem2Axi_io_dataIO_ready),
    .io_outAxi_wa_ready(mem2Axi_io_outAxi_wa_ready),
    .io_outAxi_wa_valid(mem2Axi_io_outAxi_wa_valid),
    .io_outAxi_wa_bits_id(mem2Axi_io_outAxi_wa_bits_id),
    .io_outAxi_wa_bits_addr(mem2Axi_io_outAxi_wa_bits_addr),
    .io_outAxi_wa_bits_len(mem2Axi_io_outAxi_wa_bits_len),
    .io_outAxi_wa_bits_size(mem2Axi_io_outAxi_wa_bits_size),
    .io_outAxi_wa_bits_burst(mem2Axi_io_outAxi_wa_bits_burst),
    .io_outAxi_wd_ready(mem2Axi_io_outAxi_wd_ready),
    .io_outAxi_wd_valid(mem2Axi_io_outAxi_wd_valid),
    .io_outAxi_wd_bits_data(mem2Axi_io_outAxi_wd_bits_data),
    .io_outAxi_wd_bits_strb(mem2Axi_io_outAxi_wd_bits_strb),
    .io_outAxi_wd_bits_last(mem2Axi_io_outAxi_wd_bits_last),
    .io_outAxi_wr_ready(mem2Axi_io_outAxi_wr_ready),
    .io_outAxi_wr_valid(mem2Axi_io_outAxi_wr_valid),
    .io_outAxi_wr_bits_id(mem2Axi_io_outAxi_wr_bits_id),
    .io_outAxi_wr_bits_resp(mem2Axi_io_outAxi_wr_bits_resp),
    .io_outAxi_ra_ready(mem2Axi_io_outAxi_ra_ready),
    .io_outAxi_ra_valid(mem2Axi_io_outAxi_ra_valid),
    .io_outAxi_ra_bits_id(mem2Axi_io_outAxi_ra_bits_id),
    .io_outAxi_ra_bits_addr(mem2Axi_io_outAxi_ra_bits_addr),
    .io_outAxi_ra_bits_len(mem2Axi_io_outAxi_ra_bits_len),
    .io_outAxi_ra_bits_size(mem2Axi_io_outAxi_ra_bits_size),
    .io_outAxi_ra_bits_burst(mem2Axi_io_outAxi_ra_bits_burst),
    .io_outAxi_rd_ready(mem2Axi_io_outAxi_rd_ready),
    .io_outAxi_rd_valid(mem2Axi_io_outAxi_rd_valid),
    .io_outAxi_rd_bits_id(mem2Axi_io_outAxi_rd_bits_id),
    .io_outAxi_rd_bits_data(mem2Axi_io_outAxi_rd_bits_data),
    .io_outAxi_rd_bits_resp(mem2Axi_io_outAxi_rd_bits_resp),
    .io_outAxi_rd_bits_last(mem2Axi_io_outAxi_rd_bits_last)
  );
  ysyx_210539_ToAXI flash2Axi ( // @[cpu.scala 85:29]
    .clock(flash2Axi_clock),
    .reset(flash2Axi_reset),
    .io_dataIO_addr(flash2Axi_io_dataIO_addr),
    .io_dataIO_rdata(flash2Axi_io_dataIO_rdata),
    .io_dataIO_rvalid(flash2Axi_io_dataIO_rvalid),
    .io_dataIO_wdata(flash2Axi_io_dataIO_wdata),
    .io_dataIO_dc_mode(flash2Axi_io_dataIO_dc_mode),
    .io_dataIO_ready(flash2Axi_io_dataIO_ready),
    .io_outAxi_wa_ready(flash2Axi_io_outAxi_wa_ready),
    .io_outAxi_wa_valid(flash2Axi_io_outAxi_wa_valid),
    .io_outAxi_wa_bits_id(flash2Axi_io_outAxi_wa_bits_id),
    .io_outAxi_wa_bits_addr(flash2Axi_io_outAxi_wa_bits_addr),
    .io_outAxi_wa_bits_len(flash2Axi_io_outAxi_wa_bits_len),
    .io_outAxi_wa_bits_size(flash2Axi_io_outAxi_wa_bits_size),
    .io_outAxi_wa_bits_burst(flash2Axi_io_outAxi_wa_bits_burst),
    .io_outAxi_wd_ready(flash2Axi_io_outAxi_wd_ready),
    .io_outAxi_wd_valid(flash2Axi_io_outAxi_wd_valid),
    .io_outAxi_wd_bits_data(flash2Axi_io_outAxi_wd_bits_data),
    .io_outAxi_wd_bits_strb(flash2Axi_io_outAxi_wd_bits_strb),
    .io_outAxi_wd_bits_last(flash2Axi_io_outAxi_wd_bits_last),
    .io_outAxi_wr_ready(flash2Axi_io_outAxi_wr_ready),
    .io_outAxi_wr_valid(flash2Axi_io_outAxi_wr_valid),
    .io_outAxi_wr_bits_id(flash2Axi_io_outAxi_wr_bits_id),
    .io_outAxi_wr_bits_resp(flash2Axi_io_outAxi_wr_bits_resp),
    .io_outAxi_ra_ready(flash2Axi_io_outAxi_ra_ready),
    .io_outAxi_ra_valid(flash2Axi_io_outAxi_ra_valid),
    .io_outAxi_ra_bits_id(flash2Axi_io_outAxi_ra_bits_id),
    .io_outAxi_ra_bits_addr(flash2Axi_io_outAxi_ra_bits_addr),
    .io_outAxi_ra_bits_len(flash2Axi_io_outAxi_ra_bits_len),
    .io_outAxi_ra_bits_size(flash2Axi_io_outAxi_ra_bits_size),
    .io_outAxi_ra_bits_burst(flash2Axi_io_outAxi_ra_bits_burst),
    .io_outAxi_rd_ready(flash2Axi_io_outAxi_rd_ready),
    .io_outAxi_rd_valid(flash2Axi_io_outAxi_rd_valid),
    .io_outAxi_rd_bits_id(flash2Axi_io_outAxi_rd_bits_id),
    .io_outAxi_rd_bits_data(flash2Axi_io_outAxi_rd_bits_data),
    .io_outAxi_rd_bits_resp(flash2Axi_io_outAxi_rd_bits_resp),
    .io_outAxi_rd_bits_last(flash2Axi_io_outAxi_rd_bits_last)
  );
  ysyx_210539_CrossBar crossBar ( // @[cpu.scala 87:29]
    .clock(crossBar_clock),
    .reset(crossBar_reset),
    .io_icAxi_ra_ready(crossBar_io_icAxi_ra_ready),
    .io_icAxi_ra_valid(crossBar_io_icAxi_ra_valid),
    .io_icAxi_ra_bits_addr(crossBar_io_icAxi_ra_bits_addr),
    .io_icAxi_rd_valid(crossBar_io_icAxi_rd_valid),
    .io_icAxi_rd_bits_data(crossBar_io_icAxi_rd_bits_data),
    .io_icAxi_rd_bits_last(crossBar_io_icAxi_rd_bits_last),
    .io_flashAxi_wa_ready(crossBar_io_flashAxi_wa_ready),
    .io_flashAxi_wa_valid(crossBar_io_flashAxi_wa_valid),
    .io_flashAxi_wa_bits_id(crossBar_io_flashAxi_wa_bits_id),
    .io_flashAxi_wa_bits_addr(crossBar_io_flashAxi_wa_bits_addr),
    .io_flashAxi_wa_bits_len(crossBar_io_flashAxi_wa_bits_len),
    .io_flashAxi_wa_bits_size(crossBar_io_flashAxi_wa_bits_size),
    .io_flashAxi_wa_bits_burst(crossBar_io_flashAxi_wa_bits_burst),
    .io_flashAxi_wd_ready(crossBar_io_flashAxi_wd_ready),
    .io_flashAxi_wd_valid(crossBar_io_flashAxi_wd_valid),
    .io_flashAxi_wd_bits_data(crossBar_io_flashAxi_wd_bits_data),
    .io_flashAxi_wd_bits_strb(crossBar_io_flashAxi_wd_bits_strb),
    .io_flashAxi_wd_bits_last(crossBar_io_flashAxi_wd_bits_last),
    .io_flashAxi_wr_ready(crossBar_io_flashAxi_wr_ready),
    .io_flashAxi_wr_valid(crossBar_io_flashAxi_wr_valid),
    .io_flashAxi_wr_bits_id(crossBar_io_flashAxi_wr_bits_id),
    .io_flashAxi_wr_bits_resp(crossBar_io_flashAxi_wr_bits_resp),
    .io_flashAxi_ra_ready(crossBar_io_flashAxi_ra_ready),
    .io_flashAxi_ra_valid(crossBar_io_flashAxi_ra_valid),
    .io_flashAxi_ra_bits_id(crossBar_io_flashAxi_ra_bits_id),
    .io_flashAxi_ra_bits_addr(crossBar_io_flashAxi_ra_bits_addr),
    .io_flashAxi_ra_bits_len(crossBar_io_flashAxi_ra_bits_len),
    .io_flashAxi_ra_bits_size(crossBar_io_flashAxi_ra_bits_size),
    .io_flashAxi_ra_bits_burst(crossBar_io_flashAxi_ra_bits_burst),
    .io_flashAxi_rd_ready(crossBar_io_flashAxi_rd_ready),
    .io_flashAxi_rd_valid(crossBar_io_flashAxi_rd_valid),
    .io_flashAxi_rd_bits_id(crossBar_io_flashAxi_rd_bits_id),
    .io_flashAxi_rd_bits_data(crossBar_io_flashAxi_rd_bits_data),
    .io_flashAxi_rd_bits_resp(crossBar_io_flashAxi_rd_bits_resp),
    .io_flashAxi_rd_bits_last(crossBar_io_flashAxi_rd_bits_last),
    .io_memAxi_wa_ready(crossBar_io_memAxi_wa_ready),
    .io_memAxi_wa_valid(crossBar_io_memAxi_wa_valid),
    .io_memAxi_wa_bits_addr(crossBar_io_memAxi_wa_bits_addr),
    .io_memAxi_wd_ready(crossBar_io_memAxi_wd_ready),
    .io_memAxi_wd_valid(crossBar_io_memAxi_wd_valid),
    .io_memAxi_wd_bits_data(crossBar_io_memAxi_wd_bits_data),
    .io_memAxi_wd_bits_last(crossBar_io_memAxi_wd_bits_last),
    .io_memAxi_ra_ready(crossBar_io_memAxi_ra_ready),
    .io_memAxi_ra_valid(crossBar_io_memAxi_ra_valid),
    .io_memAxi_ra_bits_addr(crossBar_io_memAxi_ra_bits_addr),
    .io_memAxi_rd_valid(crossBar_io_memAxi_rd_valid),
    .io_memAxi_rd_bits_data(crossBar_io_memAxi_rd_bits_data),
    .io_memAxi_rd_bits_last(crossBar_io_memAxi_rd_bits_last),
    .io_mmioAxi_wa_ready(crossBar_io_mmioAxi_wa_ready),
    .io_mmioAxi_wa_valid(crossBar_io_mmioAxi_wa_valid),
    .io_mmioAxi_wa_bits_id(crossBar_io_mmioAxi_wa_bits_id),
    .io_mmioAxi_wa_bits_addr(crossBar_io_mmioAxi_wa_bits_addr),
    .io_mmioAxi_wa_bits_len(crossBar_io_mmioAxi_wa_bits_len),
    .io_mmioAxi_wa_bits_size(crossBar_io_mmioAxi_wa_bits_size),
    .io_mmioAxi_wa_bits_burst(crossBar_io_mmioAxi_wa_bits_burst),
    .io_mmioAxi_wd_ready(crossBar_io_mmioAxi_wd_ready),
    .io_mmioAxi_wd_valid(crossBar_io_mmioAxi_wd_valid),
    .io_mmioAxi_wd_bits_data(crossBar_io_mmioAxi_wd_bits_data),
    .io_mmioAxi_wd_bits_strb(crossBar_io_mmioAxi_wd_bits_strb),
    .io_mmioAxi_wd_bits_last(crossBar_io_mmioAxi_wd_bits_last),
    .io_mmioAxi_wr_ready(crossBar_io_mmioAxi_wr_ready),
    .io_mmioAxi_wr_valid(crossBar_io_mmioAxi_wr_valid),
    .io_mmioAxi_wr_bits_id(crossBar_io_mmioAxi_wr_bits_id),
    .io_mmioAxi_wr_bits_resp(crossBar_io_mmioAxi_wr_bits_resp),
    .io_mmioAxi_ra_ready(crossBar_io_mmioAxi_ra_ready),
    .io_mmioAxi_ra_valid(crossBar_io_mmioAxi_ra_valid),
    .io_mmioAxi_ra_bits_id(crossBar_io_mmioAxi_ra_bits_id),
    .io_mmioAxi_ra_bits_addr(crossBar_io_mmioAxi_ra_bits_addr),
    .io_mmioAxi_ra_bits_len(crossBar_io_mmioAxi_ra_bits_len),
    .io_mmioAxi_ra_bits_size(crossBar_io_mmioAxi_ra_bits_size),
    .io_mmioAxi_ra_bits_burst(crossBar_io_mmioAxi_ra_bits_burst),
    .io_mmioAxi_rd_ready(crossBar_io_mmioAxi_rd_ready),
    .io_mmioAxi_rd_valid(crossBar_io_mmioAxi_rd_valid),
    .io_mmioAxi_rd_bits_id(crossBar_io_mmioAxi_rd_bits_id),
    .io_mmioAxi_rd_bits_data(crossBar_io_mmioAxi_rd_bits_data),
    .io_mmioAxi_rd_bits_resp(crossBar_io_mmioAxi_rd_bits_resp),
    .io_mmioAxi_rd_bits_last(crossBar_io_mmioAxi_rd_bits_last),
    .io_outAxi_wa_ready(crossBar_io_outAxi_wa_ready),
    .io_outAxi_wa_valid(crossBar_io_outAxi_wa_valid),
    .io_outAxi_wa_bits_id(crossBar_io_outAxi_wa_bits_id),
    .io_outAxi_wa_bits_addr(crossBar_io_outAxi_wa_bits_addr),
    .io_outAxi_wa_bits_len(crossBar_io_outAxi_wa_bits_len),
    .io_outAxi_wa_bits_size(crossBar_io_outAxi_wa_bits_size),
    .io_outAxi_wa_bits_burst(crossBar_io_outAxi_wa_bits_burst),
    .io_outAxi_wd_ready(crossBar_io_outAxi_wd_ready),
    .io_outAxi_wd_valid(crossBar_io_outAxi_wd_valid),
    .io_outAxi_wd_bits_data(crossBar_io_outAxi_wd_bits_data),
    .io_outAxi_wd_bits_strb(crossBar_io_outAxi_wd_bits_strb),
    .io_outAxi_wd_bits_last(crossBar_io_outAxi_wd_bits_last),
    .io_outAxi_wr_ready(crossBar_io_outAxi_wr_ready),
    .io_outAxi_wr_valid(crossBar_io_outAxi_wr_valid),
    .io_outAxi_wr_bits_id(crossBar_io_outAxi_wr_bits_id),
    .io_outAxi_wr_bits_resp(crossBar_io_outAxi_wr_bits_resp),
    .io_outAxi_ra_ready(crossBar_io_outAxi_ra_ready),
    .io_outAxi_ra_valid(crossBar_io_outAxi_ra_valid),
    .io_outAxi_ra_bits_id(crossBar_io_outAxi_ra_bits_id),
    .io_outAxi_ra_bits_addr(crossBar_io_outAxi_ra_bits_addr),
    .io_outAxi_ra_bits_len(crossBar_io_outAxi_ra_bits_len),
    .io_outAxi_ra_bits_size(crossBar_io_outAxi_ra_bits_size),
    .io_outAxi_ra_bits_burst(crossBar_io_outAxi_ra_bits_burst),
    .io_outAxi_rd_ready(crossBar_io_outAxi_rd_ready),
    .io_outAxi_rd_valid(crossBar_io_outAxi_rd_valid),
    .io_outAxi_rd_bits_id(crossBar_io_outAxi_rd_bits_id),
    .io_outAxi_rd_bits_data(crossBar_io_outAxi_rd_bits_data),
    .io_outAxi_rd_bits_resp(crossBar_io_outAxi_rd_bits_resp),
    .io_outAxi_rd_bits_last(crossBar_io_outAxi_rd_bits_last),
    .io_selectMem(crossBar_io_selectMem)
  );
  ysyx_210539_FetchCrossBar fetchCrossbar ( // @[cpu.scala 88:31]
    .clock(fetchCrossbar_clock),
    .reset(fetchCrossbar_reset),
    .io_instIO_addr(fetchCrossbar_io_instIO_addr),
    .io_instIO_inst(fetchCrossbar_io_instIO_inst),
    .io_instIO_arvalid(fetchCrossbar_io_instIO_arvalid),
    .io_instIO_rvalid(fetchCrossbar_io_instIO_rvalid),
    .io_icRead_addr(fetchCrossbar_io_icRead_addr),
    .io_icRead_inst(fetchCrossbar_io_icRead_inst),
    .io_icRead_arvalid(fetchCrossbar_io_icRead_arvalid),
    .io_icRead_rvalid(fetchCrossbar_io_icRead_rvalid),
    .io_flashRead_addr(fetchCrossbar_io_flashRead_addr),
    .io_flashRead_rdata(fetchCrossbar_io_flashRead_rdata),
    .io_flashRead_rvalid(fetchCrossbar_io_flashRead_rvalid),
    .io_flashRead_dc_mode(fetchCrossbar_io_flashRead_dc_mode)
  );
  ysyx_210539_Splite64to32 split64to32 ( // @[cpu.scala 89:29]
    .clock(split64to32_clock),
    .reset(split64to32_reset),
    .io_data_in_addr(split64to32_io_data_in_addr),
    .io_data_in_rdata(split64to32_io_data_in_rdata),
    .io_data_in_rvalid(split64to32_io_data_in_rvalid),
    .io_data_in_dc_mode(split64to32_io_data_in_dc_mode),
    .io_data_out_addr(split64to32_io_data_out_addr),
    .io_data_out_rdata(split64to32_io_data_out_rdata),
    .io_data_out_rvalid(split64to32_io_data_out_rvalid),
    .io_data_out_dc_mode(split64to32_io_data_out_dc_mode),
    .io_data_out_ready(split64to32_io_data_out_ready)
  );
  ysyx_210539_MemCrossBar memCrossbar ( // @[cpu.scala 90:29]
    .clock(memCrossbar_clock),
    .reset(memCrossbar_reset),
    .io_dataRW_addr(memCrossbar_io_dataRW_addr),
    .io_dataRW_rdata(memCrossbar_io_dataRW_rdata),
    .io_dataRW_rvalid(memCrossbar_io_dataRW_rvalid),
    .io_dataRW_wdata(memCrossbar_io_dataRW_wdata),
    .io_dataRW_dc_mode(memCrossbar_io_dataRW_dc_mode),
    .io_dataRW_amo(memCrossbar_io_dataRW_amo),
    .io_dataRW_ready(memCrossbar_io_dataRW_ready),
    .io_mmio_addr(memCrossbar_io_mmio_addr),
    .io_mmio_rdata(memCrossbar_io_mmio_rdata),
    .io_mmio_rvalid(memCrossbar_io_mmio_rvalid),
    .io_mmio_wdata(memCrossbar_io_mmio_wdata),
    .io_mmio_dc_mode(memCrossbar_io_mmio_dc_mode),
    .io_mmio_ready(memCrossbar_io_mmio_ready),
    .io_dcRW_addr(memCrossbar_io_dcRW_addr),
    .io_dcRW_rdata(memCrossbar_io_dcRW_rdata),
    .io_dcRW_rvalid(memCrossbar_io_dcRW_rvalid),
    .io_dcRW_wdata(memCrossbar_io_dcRW_wdata),
    .io_dcRW_dc_mode(memCrossbar_io_dcRW_dc_mode),
    .io_dcRW_amo(memCrossbar_io_dcRW_amo),
    .io_dcRW_ready(memCrossbar_io_dcRW_ready),
    .io_clintIO_addr(memCrossbar_io_clintIO_addr),
    .io_clintIO_rdata(memCrossbar_io_clintIO_rdata),
    .io_clintIO_wdata(memCrossbar_io_clintIO_wdata),
    .io_clintIO_wvalid(memCrossbar_io_clintIO_wvalid),
    .io_plicIO_addr(memCrossbar_io_plicIO_addr),
    .io_plicIO_rdata(memCrossbar_io_plicIO_rdata),
    .io_plicIO_wdata(memCrossbar_io_plicIO_wdata),
    .io_plicIO_wvalid(memCrossbar_io_plicIO_wvalid),
    .io_plicIO_arvalid(memCrossbar_io_plicIO_arvalid)
  );
  ysyx_210539_TLB tlb_if ( // @[cpu.scala 91:30]
    .clock(tlb_if_clock),
    .reset(tlb_if_reset),
    .io_va2pa_vaddr(tlb_if_io_va2pa_vaddr),
    .io_va2pa_vvalid(tlb_if_io_va2pa_vvalid),
    .io_va2pa_ready(tlb_if_io_va2pa_ready),
    .io_va2pa_paddr(tlb_if_io_va2pa_paddr),
    .io_va2pa_pvalid(tlb_if_io_va2pa_pvalid),
    .io_va2pa_tlb_excep_cause(tlb_if_io_va2pa_tlb_excep_cause),
    .io_va2pa_tlb_excep_tval(tlb_if_io_va2pa_tlb_excep_tval),
    .io_va2pa_tlb_excep_en(tlb_if_io_va2pa_tlb_excep_en),
    .io_mmuState_priv(tlb_if_io_mmuState_priv),
    .io_mmuState_mstatus(tlb_if_io_mmuState_mstatus),
    .io_mmuState_satp(tlb_if_io_mmuState_satp),
    .io_flush(tlb_if_io_flush),
    .io_dcacheRW_addr(tlb_if_io_dcacheRW_addr),
    .io_dcacheRW_rdata(tlb_if_io_dcacheRW_rdata),
    .io_dcacheRW_rvalid(tlb_if_io_dcacheRW_rvalid),
    .io_dcacheRW_wdata(tlb_if_io_dcacheRW_wdata),
    .io_dcacheRW_dc_mode(tlb_if_io_dcacheRW_dc_mode),
    .io_dcacheRW_ready(tlb_if_io_dcacheRW_ready)
  );
  ysyx_210539_TLB_1 tlb_mem ( // @[cpu.scala 92:30]
    .clock(tlb_mem_clock),
    .reset(tlb_mem_reset),
    .io_va2pa_vaddr(tlb_mem_io_va2pa_vaddr),
    .io_va2pa_vvalid(tlb_mem_io_va2pa_vvalid),
    .io_va2pa_m_type(tlb_mem_io_va2pa_m_type),
    .io_va2pa_ready(tlb_mem_io_va2pa_ready),
    .io_va2pa_paddr(tlb_mem_io_va2pa_paddr),
    .io_va2pa_pvalid(tlb_mem_io_va2pa_pvalid),
    .io_va2pa_tlb_excep_cause(tlb_mem_io_va2pa_tlb_excep_cause),
    .io_va2pa_tlb_excep_tval(tlb_mem_io_va2pa_tlb_excep_tval),
    .io_va2pa_tlb_excep_en(tlb_mem_io_va2pa_tlb_excep_en),
    .io_mmuState_priv(tlb_mem_io_mmuState_priv),
    .io_mmuState_mstatus(tlb_mem_io_mmuState_mstatus),
    .io_mmuState_satp(tlb_mem_io_mmuState_satp),
    .io_flush(tlb_mem_io_flush),
    .io_dcacheRW_addr(tlb_mem_io_dcacheRW_addr),
    .io_dcacheRW_rdata(tlb_mem_io_dcacheRW_rdata),
    .io_dcacheRW_rvalid(tlb_mem_io_dcacheRW_rvalid),
    .io_dcacheRW_wdata(tlb_mem_io_dcacheRW_wdata),
    .io_dcacheRW_dc_mode(tlb_mem_io_dcacheRW_dc_mode),
    .io_dcacheRW_ready(tlb_mem_io_dcacheRW_ready)
  );
  ysyx_210539_DcacheSelector dcSelector ( // @[cpu.scala 93:29]
    .clock(dcSelector_clock),
    .reset(dcSelector_reset),
    .io_tlb_if2dc_addr(dcSelector_io_tlb_if2dc_addr),
    .io_tlb_if2dc_rdata(dcSelector_io_tlb_if2dc_rdata),
    .io_tlb_if2dc_rvalid(dcSelector_io_tlb_if2dc_rvalid),
    .io_tlb_if2dc_wdata(dcSelector_io_tlb_if2dc_wdata),
    .io_tlb_if2dc_dc_mode(dcSelector_io_tlb_if2dc_dc_mode),
    .io_tlb_if2dc_ready(dcSelector_io_tlb_if2dc_ready),
    .io_tlb_mem2dc_addr(dcSelector_io_tlb_mem2dc_addr),
    .io_tlb_mem2dc_rdata(dcSelector_io_tlb_mem2dc_rdata),
    .io_tlb_mem2dc_rvalid(dcSelector_io_tlb_mem2dc_rvalid),
    .io_tlb_mem2dc_wdata(dcSelector_io_tlb_mem2dc_wdata),
    .io_tlb_mem2dc_dc_mode(dcSelector_io_tlb_mem2dc_dc_mode),
    .io_tlb_mem2dc_ready(dcSelector_io_tlb_mem2dc_ready),
    .io_mem2dc_addr(dcSelector_io_mem2dc_addr),
    .io_mem2dc_rdata(dcSelector_io_mem2dc_rdata),
    .io_mem2dc_rvalid(dcSelector_io_mem2dc_rvalid),
    .io_mem2dc_wdata(dcSelector_io_mem2dc_wdata),
    .io_mem2dc_dc_mode(dcSelector_io_mem2dc_dc_mode),
    .io_mem2dc_amo(dcSelector_io_mem2dc_amo),
    .io_mem2dc_ready(dcSelector_io_mem2dc_ready),
    .io_dma2dc_addr(dcSelector_io_dma2dc_addr),
    .io_dma2dc_rdata(dcSelector_io_dma2dc_rdata),
    .io_dma2dc_rvalid(dcSelector_io_dma2dc_rvalid),
    .io_dma2dc_wdata(dcSelector_io_dma2dc_wdata),
    .io_dma2dc_dc_mode(dcSelector_io_dma2dc_dc_mode),
    .io_dma2dc_ready(dcSelector_io_dma2dc_ready),
    .io_select_addr(dcSelector_io_select_addr),
    .io_select_rdata(dcSelector_io_select_rdata),
    .io_select_rvalid(dcSelector_io_select_rvalid),
    .io_select_wdata(dcSelector_io_select_wdata),
    .io_select_dc_mode(dcSelector_io_select_dc_mode),
    .io_select_amo(dcSelector_io_select_amo),
    .io_select_ready(dcSelector_io_select_ready)
  );
  ysyx_210539_CLINT clint ( // @[cpu.scala 94:29]
    .clock(clint_clock),
    .reset(clint_reset),
    .io_rw_addr(clint_io_rw_addr),
    .io_rw_rdata(clint_io_rw_rdata),
    .io_rw_wdata(clint_io_rw_wdata),
    .io_rw_wvalid(clint_io_rw_wvalid),
    .io_intr_raise(clint_io_intr_raise),
    .io_intr_clear(clint_io_intr_clear),
    .io_intr_msip_raise(clint_io_intr_msip_raise),
    .io_intr_msip_clear(clint_io_intr_msip_clear)
  );
  ysyx_210539_Plic plic ( // @[cpu.scala 95:29]
    .clock(plic_clock),
    .reset(plic_reset),
    .io_intr_in1(plic_io_intr_in1),
    .io_intr_out_m_raise(plic_io_intr_out_m_raise),
    .io_intr_out_m_clear(plic_io_intr_out_m_clear),
    .io_intr_out_s_raise(plic_io_intr_out_s_raise),
    .io_intr_out_s_clear(plic_io_intr_out_s_clear),
    .io_rw_addr(plic_io_rw_addr),
    .io_rw_rdata(plic_io_rw_rdata),
    .io_rw_wdata(plic_io_rw_wdata),
    .io_rw_wvalid(plic_io_rw_wvalid),
    .io_rw_arvalid(plic_io_rw_arvalid)
  );
  ysyx_210539_DmaBridge dmaBridge ( // @[cpu.scala 96:29]
    .clock(dmaBridge_clock),
    .reset(dmaBridge_reset),
    .io_dmaAxi_awready(dmaBridge_io_dmaAxi_awready),
    .io_dmaAxi_awvalid(dmaBridge_io_dmaAxi_awvalid),
    .io_dmaAxi_awaddr(dmaBridge_io_dmaAxi_awaddr),
    .io_dmaAxi_awid(dmaBridge_io_dmaAxi_awid),
    .io_dmaAxi_awlen(dmaBridge_io_dmaAxi_awlen),
    .io_dmaAxi_awsize(dmaBridge_io_dmaAxi_awsize),
    .io_dmaAxi_wready(dmaBridge_io_dmaAxi_wready),
    .io_dmaAxi_wvalid(dmaBridge_io_dmaAxi_wvalid),
    .io_dmaAxi_wdata(dmaBridge_io_dmaAxi_wdata),
    .io_dmaAxi_wstrb(dmaBridge_io_dmaAxi_wstrb),
    .io_dmaAxi_bready(dmaBridge_io_dmaAxi_bready),
    .io_dmaAxi_bvalid(dmaBridge_io_dmaAxi_bvalid),
    .io_dmaAxi_bid(dmaBridge_io_dmaAxi_bid),
    .io_dmaAxi_arready(dmaBridge_io_dmaAxi_arready),
    .io_dmaAxi_arvalid(dmaBridge_io_dmaAxi_arvalid),
    .io_dmaAxi_araddr(dmaBridge_io_dmaAxi_araddr),
    .io_dmaAxi_arid(dmaBridge_io_dmaAxi_arid),
    .io_dmaAxi_arlen(dmaBridge_io_dmaAxi_arlen),
    .io_dmaAxi_arsize(dmaBridge_io_dmaAxi_arsize),
    .io_dmaAxi_rready(dmaBridge_io_dmaAxi_rready),
    .io_dmaAxi_rvalid(dmaBridge_io_dmaAxi_rvalid),
    .io_dmaAxi_rdata(dmaBridge_io_dmaAxi_rdata),
    .io_dmaAxi_rlast(dmaBridge_io_dmaAxi_rlast),
    .io_dmaAxi_rid(dmaBridge_io_dmaAxi_rid),
    .io_dcRW_addr(dmaBridge_io_dcRW_addr),
    .io_dcRW_rdata(dmaBridge_io_dcRW_rdata),
    .io_dcRW_rvalid(dmaBridge_io_dcRW_rvalid),
    .io_dcRW_wdata(dmaBridge_io_dcRW_wdata),
    .io_dcRW_dc_mode(dmaBridge_io_dcRW_dc_mode),
    .io_dcRW_ready(dmaBridge_io_dcRW_ready)
  );
  assign io_master_awvalid = crossBar_io_outAxi_wa_valid; // @[cpu.scala 173:23]
  assign io_master_awaddr = crossBar_io_outAxi_wa_bits_addr; // @[cpu.scala 174:23]
  assign io_master_awid = crossBar_io_outAxi_wa_bits_id; // @[cpu.scala 175:23]
  assign io_master_awlen = crossBar_io_outAxi_wa_bits_len; // @[cpu.scala 176:23]
  assign io_master_awsize = crossBar_io_outAxi_wa_bits_size; // @[cpu.scala 177:23]
  assign io_master_awburst = crossBar_io_outAxi_wa_bits_burst; // @[cpu.scala 178:23]
  assign io_master_wvalid = crossBar_io_outAxi_wd_valid; // @[cpu.scala 181:23]
  assign io_master_wdata = crossBar_io_outAxi_wd_bits_data; // @[cpu.scala 182:23]
  assign io_master_wstrb = crossBar_io_outAxi_wd_bits_strb; // @[cpu.scala 183:23]
  assign io_master_wlast = crossBar_io_outAxi_wd_bits_last; // @[cpu.scala 184:23]
  assign io_master_bready = crossBar_io_outAxi_wr_ready; // @[cpu.scala 186:23]
  assign io_master_arvalid = crossBar_io_outAxi_ra_valid; // @[cpu.scala 192:23]
  assign io_master_araddr = crossBar_io_outAxi_ra_bits_addr; // @[cpu.scala 193:23]
  assign io_master_arid = crossBar_io_outAxi_ra_bits_id; // @[cpu.scala 194:23]
  assign io_master_arlen = crossBar_io_outAxi_ra_bits_len; // @[cpu.scala 195:23]
  assign io_master_arsize = crossBar_io_outAxi_ra_bits_size; // @[cpu.scala 196:23]
  assign io_master_arburst = crossBar_io_outAxi_ra_bits_burst; // @[cpu.scala 197:23]
  assign io_master_rready = crossBar_io_outAxi_rd_ready; // @[cpu.scala 199:23]
  assign io_slave_awready = dmaBridge_io_dmaAxi_awready; // @[cpu.scala 160:14]
  assign io_slave_wready = dmaBridge_io_dmaAxi_wready; // @[cpu.scala 160:14]
  assign io_slave_bvalid = dmaBridge_io_dmaAxi_bvalid; // @[cpu.scala 160:14]
  assign io_slave_bresp = 2'h0; // @[cpu.scala 160:14]
  assign io_slave_bid = dmaBridge_io_dmaAxi_bid; // @[cpu.scala 160:14]
  assign io_slave_arready = dmaBridge_io_dmaAxi_arready; // @[cpu.scala 160:14]
  assign io_slave_rvalid = dmaBridge_io_dmaAxi_rvalid; // @[cpu.scala 160:14]
  assign io_slave_rresp = 2'h0; // @[cpu.scala 160:14]
  assign io_slave_rdata = dmaBridge_io_dmaAxi_rdata; // @[cpu.scala 160:14]
  assign io_slave_rlast = dmaBridge_io_dmaAxi_rlast; // @[cpu.scala 160:14]
  assign io_slave_rid = dmaBridge_io_dmaAxi_rid; // @[cpu.scala 160:14]
  assign io_sram0_addr = icache_io_ic2sr0_addr; // @[cpu.scala 163:22]
  assign io_sram0_cen = icache_io_ic2sr0_cen; // @[cpu.scala 163:22]
  assign io_sram0_wen = icache_io_ic2sr0_wen; // @[cpu.scala 163:22]
  assign io_sram0_wmask = 128'h0; // @[cpu.scala 163:22]
  assign io_sram0_wdata = icache_io_ic2sr0_wdata; // @[cpu.scala 163:22]
  assign io_sram1_addr = icache_io_ic2sr1_addr; // @[cpu.scala 164:22]
  assign io_sram1_cen = icache_io_ic2sr1_cen; // @[cpu.scala 164:22]
  assign io_sram1_wen = icache_io_ic2sr1_wen; // @[cpu.scala 164:22]
  assign io_sram1_wmask = icache_io_ic2sr1_wmask; // @[cpu.scala 164:22]
  assign io_sram1_wdata = icache_io_ic2sr1_wdata; // @[cpu.scala 164:22]
  assign io_sram2_addr = icache_io_ic2sr2_addr; // @[cpu.scala 165:22]
  assign io_sram2_cen = icache_io_ic2sr2_cen; // @[cpu.scala 165:22]
  assign io_sram2_wen = icache_io_ic2sr2_wen; // @[cpu.scala 165:22]
  assign io_sram2_wmask = icache_io_ic2sr2_wmask; // @[cpu.scala 165:22]
  assign io_sram2_wdata = icache_io_ic2sr2_wdata; // @[cpu.scala 165:22]
  assign io_sram3_addr = icache_io_ic2sr3_addr; // @[cpu.scala 166:22]
  assign io_sram3_cen = icache_io_ic2sr3_cen; // @[cpu.scala 166:22]
  assign io_sram3_wen = icache_io_ic2sr3_wen; // @[cpu.scala 166:22]
  assign io_sram3_wmask = icache_io_ic2sr3_wmask; // @[cpu.scala 166:22]
  assign io_sram3_wdata = icache_io_ic2sr3_wdata; // @[cpu.scala 166:22]
  assign io_sram4_addr = dcache_io_dc2sr0_addr; // @[cpu.scala 167:22]
  assign io_sram4_cen = dcache_io_dc2sr0_cen; // @[cpu.scala 167:22]
  assign io_sram4_wen = dcache_io_dc2sr0_wen; // @[cpu.scala 167:22]
  assign io_sram4_wmask = dcache_io_dc2sr0_wmask; // @[cpu.scala 167:22]
  assign io_sram4_wdata = dcache_io_dc2sr0_wdata; // @[cpu.scala 167:22]
  assign io_sram5_addr = dcache_io_dc2sr1_addr; // @[cpu.scala 168:22]
  assign io_sram5_cen = dcache_io_dc2sr1_cen; // @[cpu.scala 168:22]
  assign io_sram5_wen = dcache_io_dc2sr1_wen; // @[cpu.scala 168:22]
  assign io_sram5_wmask = dcache_io_dc2sr1_wmask; // @[cpu.scala 168:22]
  assign io_sram5_wdata = dcache_io_dc2sr1_wdata; // @[cpu.scala 168:22]
  assign io_sram6_addr = dcache_io_dc2sr2_addr; // @[cpu.scala 169:22]
  assign io_sram6_cen = dcache_io_dc2sr2_cen; // @[cpu.scala 169:22]
  assign io_sram6_wen = dcache_io_dc2sr2_wen; // @[cpu.scala 169:22]
  assign io_sram6_wmask = dcache_io_dc2sr2_wmask; // @[cpu.scala 169:22]
  assign io_sram6_wdata = dcache_io_dc2sr2_wdata; // @[cpu.scala 169:22]
  assign io_sram7_addr = dcache_io_dc2sr3_addr; // @[cpu.scala 170:22]
  assign io_sram7_cen = dcache_io_dc2sr3_cen; // @[cpu.scala 170:22]
  assign io_sram7_wen = dcache_io_dc2sr3_wen; // @[cpu.scala 170:22]
  assign io_sram7_wmask = dcache_io_dc2sr3_wmask; // @[cpu.scala 170:22]
  assign io_sram7_wdata = dcache_io_dc2sr3_wdata; // @[cpu.scala 170:22]
  assign fetch_clock = clock;
  assign fetch_reset = reset;
  assign fetch_io_instRead_inst = fetchCrossbar_io_instIO_inst; // @[cpu.scala 98:25]
  assign fetch_io_instRead_rvalid = fetchCrossbar_io_instIO_rvalid; // @[cpu.scala 98:25]
  assign fetch_io_va2pa_paddr = tlb_if_io_va2pa_paddr; // @[cpu.scala 99:25]
  assign fetch_io_va2pa_pvalid = tlb_if_io_va2pa_pvalid; // @[cpu.scala 99:25]
  assign fetch_io_va2pa_tlb_excep_cause = tlb_if_io_va2pa_tlb_excep_cause; // @[cpu.scala 99:25]
  assign fetch_io_va2pa_tlb_excep_tval = tlb_if_io_va2pa_tlb_excep_tval; // @[cpu.scala 99:25]
  assign fetch_io_va2pa_tlb_excep_en = tlb_if_io_va2pa_tlb_excep_en; // @[cpu.scala 99:25]
  assign fetch_io_reg2if_seq_pc = csrs_io_reg2if_seq_pc; // @[cpu.scala 100:25]
  assign fetch_io_reg2if_valid = csrs_io_reg2if_valid; // @[cpu.scala 100:25]
  assign fetch_io_wb2if_seq_pc = writeback_io_wb2if_seq_pc; // @[cpu.scala 101:25]
  assign fetch_io_wb2if_valid = writeback_io_wb2if_valid; // @[cpu.scala 101:25]
  assign fetch_io_recov = writeback_io_recov; // @[cpu.scala 105:25]
  assign fetch_io_intr_in_en = csrs_io_intr_out_en; // @[cpu.scala 102:25]
  assign fetch_io_intr_in_cause = csrs_io_intr_out_cause; // @[cpu.scala 102:25]
  assign fetch_io_branchFail_seq_pc = execute_io_ex2if_seq_pc; // @[cpu.scala 103:25]
  assign fetch_io_branchFail_valid = execute_io_ex2if_valid; // @[cpu.scala 103:25]
  assign fetch_io_if2id_drop = decode_io_if2id_drop; // @[cpu.scala 104:25]
  assign fetch_io_if2id_stall = decode_io_if2id_stall; // @[cpu.scala 104:25]
  assign fetch_io_if2id_ready = decode_io_if2id_ready; // @[cpu.scala 104:25]
  assign decode_clock = clock;
  assign decode_reset = reset;
  assign decode_io_if2id_inst = fetch_io_if2id_inst; // @[cpu.scala 104:25]
  assign decode_io_if2id_pc = fetch_io_if2id_pc; // @[cpu.scala 104:25]
  assign decode_io_if2id_excep_cause = fetch_io_if2id_excep_cause; // @[cpu.scala 104:25]
  assign decode_io_if2id_excep_tval = fetch_io_if2id_excep_tval; // @[cpu.scala 104:25]
  assign decode_io_if2id_excep_en = fetch_io_if2id_excep_en; // @[cpu.scala 104:25]
  assign decode_io_if2id_excep_pc = fetch_io_if2id_excep_pc; // @[cpu.scala 104:25]
  assign decode_io_if2id_recov = fetch_io_if2id_recov; // @[cpu.scala 104:25]
  assign decode_io_if2id_valid = fetch_io_if2id_valid; // @[cpu.scala 104:25]
  assign decode_io_id2df_drop = forwading_io_id2df_drop; // @[cpu.scala 107:25]
  assign decode_io_id2df_stall = forwading_io_id2df_stall; // @[cpu.scala 107:25]
  assign decode_io_id2df_ready = forwading_io_id2df_ready; // @[cpu.scala 107:25]
  assign decode_io_idState_priv = csrs_io_idState_priv; // @[cpu.scala 108:25]
  assign forwading_clock = clock;
  assign forwading_reset = reset;
  assign forwading_io_id2df_inst = decode_io_id2df_inst; // @[cpu.scala 107:25]
  assign forwading_io_id2df_pc = decode_io_id2df_pc; // @[cpu.scala 107:25]
  assign forwading_io_id2df_excep_cause = decode_io_id2df_excep_cause; // @[cpu.scala 107:25]
  assign forwading_io_id2df_excep_tval = decode_io_id2df_excep_tval; // @[cpu.scala 107:25]
  assign forwading_io_id2df_excep_en = decode_io_id2df_excep_en; // @[cpu.scala 107:25]
  assign forwading_io_id2df_excep_pc = decode_io_id2df_excep_pc; // @[cpu.scala 107:25]
  assign forwading_io_id2df_excep_etype = decode_io_id2df_excep_etype; // @[cpu.scala 107:25]
  assign forwading_io_id2df_ctrl_aluOp = decode_io_id2df_ctrl_aluOp; // @[cpu.scala 107:25]
  assign forwading_io_id2df_ctrl_aluWidth = decode_io_id2df_ctrl_aluWidth; // @[cpu.scala 107:25]
  assign forwading_io_id2df_ctrl_dcMode = decode_io_id2df_ctrl_dcMode; // @[cpu.scala 107:25]
  assign forwading_io_id2df_ctrl_writeRegEn = decode_io_id2df_ctrl_writeRegEn; // @[cpu.scala 107:25]
  assign forwading_io_id2df_ctrl_writeCSREn = decode_io_id2df_ctrl_writeCSREn; // @[cpu.scala 107:25]
  assign forwading_io_id2df_ctrl_brType = decode_io_id2df_ctrl_brType; // @[cpu.scala 107:25]
  assign forwading_io_id2df_rs1 = decode_io_id2df_rs1; // @[cpu.scala 107:25]
  assign forwading_io_id2df_rrs1 = decode_io_id2df_rrs1; // @[cpu.scala 107:25]
  assign forwading_io_id2df_rs1_d = decode_io_id2df_rs1_d; // @[cpu.scala 107:25]
  assign forwading_io_id2df_rs2 = decode_io_id2df_rs2; // @[cpu.scala 107:25]
  assign forwading_io_id2df_rrs2 = decode_io_id2df_rrs2; // @[cpu.scala 107:25]
  assign forwading_io_id2df_rs2_d = decode_io_id2df_rs2_d; // @[cpu.scala 107:25]
  assign forwading_io_id2df_dst = decode_io_id2df_dst; // @[cpu.scala 107:25]
  assign forwading_io_id2df_dst_d = decode_io_id2df_dst_d; // @[cpu.scala 107:25]
  assign forwading_io_id2df_jmp_type = decode_io_id2df_jmp_type; // @[cpu.scala 107:25]
  assign forwading_io_id2df_special = decode_io_id2df_special; // @[cpu.scala 107:25]
  assign forwading_io_id2df_swap = decode_io_id2df_swap; // @[cpu.scala 107:25]
  assign forwading_io_id2df_indi = decode_io_id2df_indi; // @[cpu.scala 107:25]
  assign forwading_io_id2df_recov = decode_io_id2df_recov; // @[cpu.scala 107:25]
  assign forwading_io_id2df_valid = decode_io_id2df_valid; // @[cpu.scala 107:25]
  assign forwading_io_df2rr_drop = readregs_io_df2rr_drop; // @[cpu.scala 109:25]
  assign forwading_io_df2rr_stall = readregs_io_df2rr_stall; // @[cpu.scala 109:25]
  assign forwading_io_df2rr_ready = readregs_io_df2rr_ready; // @[cpu.scala 109:25]
  assign forwading_io_d_rr_id = readregs_io_d_rr_id; // @[cpu.scala 110:25]
  assign forwading_io_d_rr_data = readregs_io_d_rr_data; // @[cpu.scala 110:25]
  assign forwading_io_d_rr_state = readregs_io_d_rr_state; // @[cpu.scala 110:25]
  assign forwading_io_d_ex_id = execute_io_d_ex_id; // @[cpu.scala 111:25]
  assign forwading_io_d_ex_data = execute_io_d_ex_data; // @[cpu.scala 111:25]
  assign forwading_io_d_ex_state = execute_io_d_ex_state; // @[cpu.scala 111:25]
  assign forwading_io_d_mem1_id = memory_io_d_mem1_id; // @[cpu.scala 112:25]
  assign forwading_io_d_mem1_data = memory_io_d_mem1_data; // @[cpu.scala 112:25]
  assign forwading_io_d_mem1_state = memory_io_d_mem1_state; // @[cpu.scala 112:25]
  assign forwading_io_d_mem2_id = memory_io_d_mem2_id; // @[cpu.scala 113:25]
  assign forwading_io_d_mem2_data = memory_io_d_mem2_data; // @[cpu.scala 113:25]
  assign forwading_io_d_mem2_state = memory_io_d_mem2_state; // @[cpu.scala 113:25]
  assign forwading_io_d_mem3_id = memory_io_d_mem3_id; // @[cpu.scala 114:25]
  assign forwading_io_d_mem3_data = memory_io_d_mem3_data; // @[cpu.scala 114:25]
  assign forwading_io_d_mem3_state = memory_io_d_mem3_state; // @[cpu.scala 114:25]
  assign readregs_clock = clock;
  assign readregs_reset = reset;
  assign readregs_io_df2rr_inst = forwading_io_df2rr_inst; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_pc = forwading_io_df2rr_pc; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_excep_cause = forwading_io_df2rr_excep_cause; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_excep_tval = forwading_io_df2rr_excep_tval; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_excep_en = forwading_io_df2rr_excep_en; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_excep_pc = forwading_io_df2rr_excep_pc; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_excep_etype = forwading_io_df2rr_excep_etype; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_ctrl_aluOp = forwading_io_df2rr_ctrl_aluOp; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_ctrl_aluWidth = forwading_io_df2rr_ctrl_aluWidth; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_ctrl_dcMode = forwading_io_df2rr_ctrl_dcMode; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_ctrl_writeRegEn = forwading_io_df2rr_ctrl_writeRegEn; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_ctrl_writeCSREn = forwading_io_df2rr_ctrl_writeCSREn; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_ctrl_brType = forwading_io_df2rr_ctrl_brType; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_rs1 = forwading_io_df2rr_rs1; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_rrs1 = forwading_io_df2rr_rrs1; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_rs1_d = forwading_io_df2rr_rs1_d; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_rs2 = forwading_io_df2rr_rs2; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_rrs2 = forwading_io_df2rr_rrs2; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_rs2_d = forwading_io_df2rr_rs2_d; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_dst = forwading_io_df2rr_dst; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_dst_d = forwading_io_df2rr_dst_d; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_jmp_type = forwading_io_df2rr_jmp_type; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_special = forwading_io_df2rr_special; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_swap = forwading_io_df2rr_swap; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_indi = forwading_io_df2rr_indi; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_recov = forwading_io_df2rr_recov; // @[cpu.scala 109:25]
  assign readregs_io_df2rr_valid = forwading_io_df2rr_valid; // @[cpu.scala 109:25]
  assign readregs_io_rr2ex_drop = execute_io_rr2ex_drop; // @[cpu.scala 115:25]
  assign readregs_io_rr2ex_stall = execute_io_rr2ex_stall; // @[cpu.scala 115:25]
  assign readregs_io_rr2ex_ready = execute_io_rr2ex_ready; // @[cpu.scala 115:25]
  assign readregs_io_rs1Read_data = regs_io_rs1_data; // @[cpu.scala 116:25]
  assign readregs_io_rs2Read_data = regs_io_rs2_data; // @[cpu.scala 117:25]
  assign readregs_io_csrRead_data = csrs_io_rs_data; // @[cpu.scala 118:25]
  assign readregs_io_csrRead_is_err = csrs_io_rs_is_err; // @[cpu.scala 118:25]
  assign execute_clock = clock;
  assign execute_reset = reset;
  assign execute_io_rr2ex_inst = readregs_io_rr2ex_inst; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_pc = readregs_io_rr2ex_pc; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_excep_cause = readregs_io_rr2ex_excep_cause; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_excep_tval = readregs_io_rr2ex_excep_tval; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_excep_en = readregs_io_rr2ex_excep_en; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_excep_pc = readregs_io_rr2ex_excep_pc; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_excep_etype = readregs_io_rr2ex_excep_etype; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_ctrl_aluOp = readregs_io_rr2ex_ctrl_aluOp; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_ctrl_aluWidth = readregs_io_rr2ex_ctrl_aluWidth; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_ctrl_dcMode = readregs_io_rr2ex_ctrl_dcMode; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_ctrl_writeRegEn = readregs_io_rr2ex_ctrl_writeRegEn; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_ctrl_writeCSREn = readregs_io_rr2ex_ctrl_writeCSREn; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_ctrl_brType = readregs_io_rr2ex_ctrl_brType; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_rs1_d = readregs_io_rr2ex_rs1_d; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_rs2 = readregs_io_rr2ex_rs2; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_rs2_d = readregs_io_rr2ex_rs2_d; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_dst = readregs_io_rr2ex_dst; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_dst_d = readregs_io_rr2ex_dst_d; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_rcsr_id = readregs_io_rr2ex_rcsr_id; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_jmp_type = readregs_io_rr2ex_jmp_type; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_special = readregs_io_rr2ex_special; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_indi = readregs_io_rr2ex_indi; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_recov = readregs_io_rr2ex_recov; // @[cpu.scala 115:25]
  assign execute_io_rr2ex_valid = readregs_io_rr2ex_valid; // @[cpu.scala 115:25]
  assign execute_io_ex2mem_drop = memory_io_ex2mem_drop; // @[cpu.scala 120:25]
  assign execute_io_ex2mem_stall = memory_io_ex2mem_stall; // @[cpu.scala 120:25]
  assign execute_io_ex2mem_ready = memory_io_ex2mem_ready; // @[cpu.scala 120:25]
  assign execute_io_updateNextPc_seq_pc = csrs_io_updateNextPc_seq_pc; // @[cpu.scala 121:29]
  assign execute_io_updateNextPc_valid = csrs_io_updateNextPc_valid; // @[cpu.scala 121:29]
  assign memory_clock = clock;
  assign memory_reset = reset;
  assign memory_io_ex2mem_inst = execute_io_ex2mem_inst; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_pc = execute_io_ex2mem_pc; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_excep_cause = execute_io_ex2mem_excep_cause; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_excep_tval = execute_io_ex2mem_excep_tval; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_excep_en = execute_io_ex2mem_excep_en; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_excep_pc = execute_io_ex2mem_excep_pc; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_excep_etype = execute_io_ex2mem_excep_etype; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_ctrl_dcMode = execute_io_ex2mem_ctrl_dcMode; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_ctrl_writeRegEn = execute_io_ex2mem_ctrl_writeRegEn; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_ctrl_writeCSREn = execute_io_ex2mem_ctrl_writeCSREn; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_mem_addr = execute_io_ex2mem_mem_addr; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_mem_data = execute_io_ex2mem_mem_data; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_csr_id = execute_io_ex2mem_csr_id; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_csr_d = execute_io_ex2mem_csr_d; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_dst = execute_io_ex2mem_dst; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_dst_d = execute_io_ex2mem_dst_d; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_rcsr_id = execute_io_ex2mem_rcsr_id; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_special = execute_io_ex2mem_special; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_indi = execute_io_ex2mem_indi; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_recov = execute_io_ex2mem_recov; // @[cpu.scala 120:25]
  assign memory_io_ex2mem_valid = execute_io_ex2mem_valid; // @[cpu.scala 120:25]
  assign memory_io_mem2rb_drop = writeback_io_mem2rb_drop; // @[cpu.scala 122:25]
  assign memory_io_mem2rb_stall = writeback_io_mem2rb_stall; // @[cpu.scala 122:25]
  assign memory_io_mem2rb_ready = writeback_io_mem2rb_ready; // @[cpu.scala 122:25]
  assign memory_io_dataRW_rdata = memCrossbar_io_dataRW_rdata; // @[cpu.scala 123:25]
  assign memory_io_dataRW_rvalid = memCrossbar_io_dataRW_rvalid; // @[cpu.scala 123:25]
  assign memory_io_dataRW_ready = memCrossbar_io_dataRW_ready; // @[cpu.scala 123:25]
  assign memory_io_va2pa_paddr = tlb_mem_io_va2pa_paddr; // @[cpu.scala 124:25]
  assign memory_io_va2pa_pvalid = tlb_mem_io_va2pa_pvalid; // @[cpu.scala 124:25]
  assign memory_io_va2pa_tlb_excep_cause = tlb_mem_io_va2pa_tlb_excep_cause; // @[cpu.scala 124:25]
  assign memory_io_va2pa_tlb_excep_tval = tlb_mem_io_va2pa_tlb_excep_tval; // @[cpu.scala 124:25]
  assign memory_io_va2pa_tlb_excep_en = tlb_mem_io_va2pa_tlb_excep_en; // @[cpu.scala 124:25]
  assign writeback_clock = clock;
  assign writeback_reset = reset;
  assign writeback_io_mem2rb_inst = memory_io_mem2rb_inst; // @[cpu.scala 122:25]
  assign writeback_io_mem2rb_pc = memory_io_mem2rb_pc; // @[cpu.scala 122:25]
  assign writeback_io_mem2rb_excep_cause = memory_io_mem2rb_excep_cause; // @[cpu.scala 122:25]
  assign writeback_io_mem2rb_excep_tval = memory_io_mem2rb_excep_tval; // @[cpu.scala 122:25]
  assign writeback_io_mem2rb_excep_en = memory_io_mem2rb_excep_en; // @[cpu.scala 122:25]
  assign writeback_io_mem2rb_excep_pc = memory_io_mem2rb_excep_pc; // @[cpu.scala 122:25]
  assign writeback_io_mem2rb_excep_etype = memory_io_mem2rb_excep_etype; // @[cpu.scala 122:25]
  assign writeback_io_mem2rb_csr_id = memory_io_mem2rb_csr_id; // @[cpu.scala 122:25]
  assign writeback_io_mem2rb_csr_d = memory_io_mem2rb_csr_d; // @[cpu.scala 122:25]
  assign writeback_io_mem2rb_csr_en = memory_io_mem2rb_csr_en; // @[cpu.scala 122:25]
  assign writeback_io_mem2rb_dst = memory_io_mem2rb_dst; // @[cpu.scala 122:25]
  assign writeback_io_mem2rb_dst_d = memory_io_mem2rb_dst_d; // @[cpu.scala 122:25]
  assign writeback_io_mem2rb_dst_en = memory_io_mem2rb_dst_en; // @[cpu.scala 122:25]
  assign writeback_io_mem2rb_rcsr_id = memory_io_mem2rb_rcsr_id; // @[cpu.scala 122:25]
  assign writeback_io_mem2rb_special = memory_io_mem2rb_special; // @[cpu.scala 122:25]
  assign writeback_io_mem2rb_is_mmio = memory_io_mem2rb_is_mmio; // @[cpu.scala 122:25]
  assign writeback_io_mem2rb_recov = memory_io_mem2rb_recov; // @[cpu.scala 122:25]
  assign writeback_io_mem2rb_valid = memory_io_mem2rb_valid; // @[cpu.scala 122:25]
  assign regs_clock = clock;
  assign regs_reset = reset;
  assign regs_io_rs1_id = readregs_io_rs1Read_id; // @[cpu.scala 116:25]
  assign regs_io_rs2_id = readregs_io_rs2Read_id; // @[cpu.scala 117:25]
  assign regs_io_dst_id = writeback_io_wReg_id; // @[cpu.scala 126:25]
  assign regs_io_dst_data = writeback_io_wReg_data; // @[cpu.scala 126:25]
  assign regs_io_dst_en = writeback_io_wReg_en; // @[cpu.scala 126:25]
  assign csrs_clock = clock;
  assign csrs_reset = reset;
  assign csrs_io_rs_id = readregs_io_csrRead_id; // @[cpu.scala 118:25]
  assign csrs_io_rd_id = writeback_io_wCsr_id; // @[cpu.scala 127:25]
  assign csrs_io_rd_data = writeback_io_wCsr_data; // @[cpu.scala 127:25]
  assign csrs_io_rd_en = writeback_io_wCsr_en; // @[cpu.scala 127:25]
  assign csrs_io_excep_cause = writeback_io_excep_cause; // @[cpu.scala 128:25]
  assign csrs_io_excep_tval = writeback_io_excep_tval; // @[cpu.scala 128:25]
  assign csrs_io_excep_en = writeback_io_excep_en; // @[cpu.scala 128:25]
  assign csrs_io_excep_pc = writeback_io_excep_pc; // @[cpu.scala 128:25]
  assign csrs_io_excep_etype = writeback_io_excep_etype; // @[cpu.scala 128:25]
  assign csrs_io_clint_raise = clint_io_intr_raise; // @[cpu.scala 129:25]
  assign csrs_io_clint_clear = clint_io_intr_clear; // @[cpu.scala 129:25]
  assign csrs_io_plic_m_raise = plic_io_intr_out_m_raise; // @[cpu.scala 156:25]
  assign csrs_io_plic_m_clear = plic_io_intr_out_m_clear; // @[cpu.scala 156:25]
  assign csrs_io_plic_s_raise = plic_io_intr_out_s_raise; // @[cpu.scala 157:25]
  assign csrs_io_plic_s_clear = plic_io_intr_out_s_clear; // @[cpu.scala 157:25]
  assign csrs_io_intr_msip_raise = clint_io_intr_msip_raise; // @[cpu.scala 130:25]
  assign csrs_io_intr_msip_clear = clint_io_intr_msip_clear; // @[cpu.scala 130:25]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_instAxi_ra_ready = crossBar_io_icAxi_ra_ready; // @[cpu.scala 149:25]
  assign icache_io_instAxi_rd_valid = crossBar_io_icAxi_rd_valid; // @[cpu.scala 149:25]
  assign icache_io_instAxi_rd_bits_data = crossBar_io_icAxi_rd_bits_data; // @[cpu.scala 149:25]
  assign icache_io_instAxi_rd_bits_last = crossBar_io_icAxi_rd_bits_last; // @[cpu.scala 149:25]
  assign icache_io_icRead_addr = fetchCrossbar_io_icRead_addr; // @[cpu.scala 137:33]
  assign icache_io_icRead_arvalid = fetchCrossbar_io_icRead_arvalid; // @[cpu.scala 137:33]
  assign icache_io_flush = writeback_io_flush_cache; // @[cpu.scala 132:25]
  assign icache_io_ic2sr0_rdata = io_sram0_rdata; // @[cpu.scala 163:22]
  assign icache_io_ic2sr1_rdata = io_sram1_rdata; // @[cpu.scala 164:22]
  assign icache_io_ic2sr2_rdata = io_sram2_rdata; // @[cpu.scala 165:22]
  assign icache_io_ic2sr3_rdata = io_sram3_rdata; // @[cpu.scala 166:22]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_dataAxi_wa_ready = crossBar_io_memAxi_wa_ready; // @[cpu.scala 150:25]
  assign dcache_io_dataAxi_wd_ready = crossBar_io_memAxi_wd_ready; // @[cpu.scala 150:25]
  assign dcache_io_dataAxi_ra_ready = crossBar_io_memAxi_ra_ready; // @[cpu.scala 150:25]
  assign dcache_io_dataAxi_rd_valid = crossBar_io_memAxi_rd_valid; // @[cpu.scala 150:25]
  assign dcache_io_dataAxi_rd_bits_data = crossBar_io_memAxi_rd_bits_data; // @[cpu.scala 150:25]
  assign dcache_io_dataAxi_rd_bits_last = crossBar_io_memAxi_rd_bits_last; // @[cpu.scala 150:25]
  assign dcache_io_dcRW_addr = dcSelector_io_select_addr; // @[cpu.scala 143:33]
  assign dcache_io_dcRW_wdata = dcSelector_io_select_wdata; // @[cpu.scala 143:33]
  assign dcache_io_dcRW_dc_mode = dcSelector_io_select_dc_mode; // @[cpu.scala 143:33]
  assign dcache_io_dcRW_amo = dcSelector_io_select_amo; // @[cpu.scala 143:33]
  assign dcache_io_flush = writeback_io_flush_cache; // @[cpu.scala 133:25]
  assign dcache_io_dc2sr0_rdata = io_sram4_rdata; // @[cpu.scala 167:22]
  assign dcache_io_dc2sr1_rdata = io_sram5_rdata; // @[cpu.scala 168:22]
  assign dcache_io_dc2sr2_rdata = io_sram6_rdata; // @[cpu.scala 169:22]
  assign dcache_io_dc2sr3_rdata = io_sram7_rdata; // @[cpu.scala 170:22]
  assign mem2Axi_clock = clock;
  assign mem2Axi_reset = reset;
  assign mem2Axi_io_dataIO_addr = memCrossbar_io_mmio_addr; // @[cpu.scala 141:33]
  assign mem2Axi_io_dataIO_wdata = memCrossbar_io_mmio_wdata; // @[cpu.scala 141:33]
  assign mem2Axi_io_dataIO_dc_mode = memCrossbar_io_mmio_dc_mode; // @[cpu.scala 141:33]
  assign mem2Axi_io_outAxi_wa_ready = crossBar_io_mmioAxi_wa_ready; // @[cpu.scala 151:25]
  assign mem2Axi_io_outAxi_wd_ready = crossBar_io_mmioAxi_wd_ready; // @[cpu.scala 151:25]
  assign mem2Axi_io_outAxi_wr_valid = crossBar_io_mmioAxi_wr_valid; // @[cpu.scala 151:25]
  assign mem2Axi_io_outAxi_wr_bits_id = crossBar_io_mmioAxi_wr_bits_id; // @[cpu.scala 151:25]
  assign mem2Axi_io_outAxi_wr_bits_resp = crossBar_io_mmioAxi_wr_bits_resp; // @[cpu.scala 151:25]
  assign mem2Axi_io_outAxi_ra_ready = crossBar_io_mmioAxi_ra_ready; // @[cpu.scala 151:25]
  assign mem2Axi_io_outAxi_rd_valid = crossBar_io_mmioAxi_rd_valid; // @[cpu.scala 151:25]
  assign mem2Axi_io_outAxi_rd_bits_id = crossBar_io_mmioAxi_rd_bits_id; // @[cpu.scala 151:25]
  assign mem2Axi_io_outAxi_rd_bits_data = crossBar_io_mmioAxi_rd_bits_data; // @[cpu.scala 151:25]
  assign mem2Axi_io_outAxi_rd_bits_resp = crossBar_io_mmioAxi_rd_bits_resp; // @[cpu.scala 151:25]
  assign mem2Axi_io_outAxi_rd_bits_last = crossBar_io_mmioAxi_rd_bits_last; // @[cpu.scala 151:25]
  assign flash2Axi_clock = clock;
  assign flash2Axi_reset = reset;
  assign flash2Axi_io_dataIO_addr = split64to32_io_data_out_addr; // @[cpu.scala 139:33]
  assign flash2Axi_io_dataIO_wdata = 64'h0; // @[cpu.scala 139:33]
  assign flash2Axi_io_dataIO_dc_mode = split64to32_io_data_out_dc_mode; // @[cpu.scala 139:33]
  assign flash2Axi_io_outAxi_wa_ready = crossBar_io_flashAxi_wa_ready; // @[cpu.scala 152:26]
  assign flash2Axi_io_outAxi_wd_ready = crossBar_io_flashAxi_wd_ready; // @[cpu.scala 152:26]
  assign flash2Axi_io_outAxi_wr_valid = crossBar_io_flashAxi_wr_valid; // @[cpu.scala 152:26]
  assign flash2Axi_io_outAxi_wr_bits_id = crossBar_io_flashAxi_wr_bits_id; // @[cpu.scala 152:26]
  assign flash2Axi_io_outAxi_wr_bits_resp = crossBar_io_flashAxi_wr_bits_resp; // @[cpu.scala 152:26]
  assign flash2Axi_io_outAxi_ra_ready = crossBar_io_flashAxi_ra_ready; // @[cpu.scala 152:26]
  assign flash2Axi_io_outAxi_rd_valid = crossBar_io_flashAxi_rd_valid; // @[cpu.scala 152:26]
  assign flash2Axi_io_outAxi_rd_bits_id = crossBar_io_flashAxi_rd_bits_id; // @[cpu.scala 152:26]
  assign flash2Axi_io_outAxi_rd_bits_data = crossBar_io_flashAxi_rd_bits_data; // @[cpu.scala 152:26]
  assign flash2Axi_io_outAxi_rd_bits_resp = crossBar_io_flashAxi_rd_bits_resp; // @[cpu.scala 152:26]
  assign flash2Axi_io_outAxi_rd_bits_last = crossBar_io_flashAxi_rd_bits_last; // @[cpu.scala 152:26]
  assign crossBar_clock = clock;
  assign crossBar_reset = reset;
  assign crossBar_io_icAxi_ra_valid = icache_io_instAxi_ra_valid; // @[cpu.scala 149:25]
  assign crossBar_io_icAxi_ra_bits_addr = icache_io_instAxi_ra_bits_addr; // @[cpu.scala 149:25]
  assign crossBar_io_flashAxi_wa_valid = flash2Axi_io_outAxi_wa_valid; // @[cpu.scala 152:26]
  assign crossBar_io_flashAxi_wa_bits_id = flash2Axi_io_outAxi_wa_bits_id; // @[cpu.scala 152:26]
  assign crossBar_io_flashAxi_wa_bits_addr = flash2Axi_io_outAxi_wa_bits_addr; // @[cpu.scala 152:26]
  assign crossBar_io_flashAxi_wa_bits_len = flash2Axi_io_outAxi_wa_bits_len; // @[cpu.scala 152:26]
  assign crossBar_io_flashAxi_wa_bits_size = flash2Axi_io_outAxi_wa_bits_size; // @[cpu.scala 152:26]
  assign crossBar_io_flashAxi_wa_bits_burst = flash2Axi_io_outAxi_wa_bits_burst; // @[cpu.scala 152:26]
  assign crossBar_io_flashAxi_wd_valid = flash2Axi_io_outAxi_wd_valid; // @[cpu.scala 152:26]
  assign crossBar_io_flashAxi_wd_bits_data = flash2Axi_io_outAxi_wd_bits_data; // @[cpu.scala 152:26]
  assign crossBar_io_flashAxi_wd_bits_strb = flash2Axi_io_outAxi_wd_bits_strb; // @[cpu.scala 152:26]
  assign crossBar_io_flashAxi_wd_bits_last = flash2Axi_io_outAxi_wd_bits_last; // @[cpu.scala 152:26]
  assign crossBar_io_flashAxi_wr_ready = flash2Axi_io_outAxi_wr_ready; // @[cpu.scala 152:26]
  assign crossBar_io_flashAxi_ra_valid = flash2Axi_io_outAxi_ra_valid; // @[cpu.scala 152:26]
  assign crossBar_io_flashAxi_ra_bits_id = flash2Axi_io_outAxi_ra_bits_id; // @[cpu.scala 152:26]
  assign crossBar_io_flashAxi_ra_bits_addr = flash2Axi_io_outAxi_ra_bits_addr; // @[cpu.scala 152:26]
  assign crossBar_io_flashAxi_ra_bits_len = flash2Axi_io_outAxi_ra_bits_len; // @[cpu.scala 152:26]
  assign crossBar_io_flashAxi_ra_bits_size = flash2Axi_io_outAxi_ra_bits_size; // @[cpu.scala 152:26]
  assign crossBar_io_flashAxi_ra_bits_burst = flash2Axi_io_outAxi_ra_bits_burst; // @[cpu.scala 152:26]
  assign crossBar_io_flashAxi_rd_ready = flash2Axi_io_outAxi_rd_ready; // @[cpu.scala 152:26]
  assign crossBar_io_memAxi_wa_valid = dcache_io_dataAxi_wa_valid; // @[cpu.scala 150:25]
  assign crossBar_io_memAxi_wa_bits_addr = dcache_io_dataAxi_wa_bits_addr; // @[cpu.scala 150:25]
  assign crossBar_io_memAxi_wd_valid = dcache_io_dataAxi_wd_valid; // @[cpu.scala 150:25]
  assign crossBar_io_memAxi_wd_bits_data = dcache_io_dataAxi_wd_bits_data; // @[cpu.scala 150:25]
  assign crossBar_io_memAxi_wd_bits_last = dcache_io_dataAxi_wd_bits_last; // @[cpu.scala 150:25]
  assign crossBar_io_memAxi_ra_valid = dcache_io_dataAxi_ra_valid; // @[cpu.scala 150:25]
  assign crossBar_io_memAxi_ra_bits_addr = dcache_io_dataAxi_ra_bits_addr; // @[cpu.scala 150:25]
  assign crossBar_io_mmioAxi_wa_valid = mem2Axi_io_outAxi_wa_valid; // @[cpu.scala 151:25]
  assign crossBar_io_mmioAxi_wa_bits_id = mem2Axi_io_outAxi_wa_bits_id; // @[cpu.scala 151:25]
  assign crossBar_io_mmioAxi_wa_bits_addr = mem2Axi_io_outAxi_wa_bits_addr; // @[cpu.scala 151:25]
  assign crossBar_io_mmioAxi_wa_bits_len = mem2Axi_io_outAxi_wa_bits_len; // @[cpu.scala 151:25]
  assign crossBar_io_mmioAxi_wa_bits_size = mem2Axi_io_outAxi_wa_bits_size; // @[cpu.scala 151:25]
  assign crossBar_io_mmioAxi_wa_bits_burst = mem2Axi_io_outAxi_wa_bits_burst; // @[cpu.scala 151:25]
  assign crossBar_io_mmioAxi_wd_valid = mem2Axi_io_outAxi_wd_valid; // @[cpu.scala 151:25]
  assign crossBar_io_mmioAxi_wd_bits_data = mem2Axi_io_outAxi_wd_bits_data; // @[cpu.scala 151:25]
  assign crossBar_io_mmioAxi_wd_bits_strb = mem2Axi_io_outAxi_wd_bits_strb; // @[cpu.scala 151:25]
  assign crossBar_io_mmioAxi_wd_bits_last = mem2Axi_io_outAxi_wd_bits_last; // @[cpu.scala 151:25]
  assign crossBar_io_mmioAxi_wr_ready = mem2Axi_io_outAxi_wr_ready; // @[cpu.scala 151:25]
  assign crossBar_io_mmioAxi_ra_valid = mem2Axi_io_outAxi_ra_valid; // @[cpu.scala 151:25]
  assign crossBar_io_mmioAxi_ra_bits_id = mem2Axi_io_outAxi_ra_bits_id; // @[cpu.scala 151:25]
  assign crossBar_io_mmioAxi_ra_bits_addr = mem2Axi_io_outAxi_ra_bits_addr; // @[cpu.scala 151:25]
  assign crossBar_io_mmioAxi_ra_bits_len = mem2Axi_io_outAxi_ra_bits_len; // @[cpu.scala 151:25]
  assign crossBar_io_mmioAxi_ra_bits_size = mem2Axi_io_outAxi_ra_bits_size; // @[cpu.scala 151:25]
  assign crossBar_io_mmioAxi_ra_bits_burst = mem2Axi_io_outAxi_ra_bits_burst; // @[cpu.scala 151:25]
  assign crossBar_io_mmioAxi_rd_ready = mem2Axi_io_outAxi_rd_ready; // @[cpu.scala 151:25]
  assign crossBar_io_outAxi_wa_ready = io_master_awready; // @[cpu.scala 172:36]
  assign crossBar_io_outAxi_wd_ready = io_master_wready; // @[cpu.scala 180:35]
  assign crossBar_io_outAxi_wr_valid = io_master_bvalid; // @[cpu.scala 187:40]
  assign crossBar_io_outAxi_wr_bits_id = io_master_bid; // @[cpu.scala 189:40]
  assign crossBar_io_outAxi_wr_bits_resp = io_master_bresp; // @[cpu.scala 188:40]
  assign crossBar_io_outAxi_ra_ready = io_master_arready; // @[cpu.scala 191:34]
  assign crossBar_io_outAxi_rd_valid = io_master_rvalid; // @[cpu.scala 200:35]
  assign crossBar_io_outAxi_rd_bits_id = io_master_rid; // @[cpu.scala 204:40]
  assign crossBar_io_outAxi_rd_bits_data = io_master_rdata; // @[cpu.scala 202:40]
  assign crossBar_io_outAxi_rd_bits_resp = io_master_rresp; // @[cpu.scala 201:40]
  assign crossBar_io_outAxi_rd_bits_last = io_master_rlast; // @[cpu.scala 203:40]
  assign crossBar_io_selectMem = dcache_io_flush_out; // @[cpu.scala 153:27]
  assign fetchCrossbar_clock = clock;
  assign fetchCrossbar_reset = reset;
  assign fetchCrossbar_io_instIO_addr = fetch_io_instRead_addr; // @[cpu.scala 98:25]
  assign fetchCrossbar_io_instIO_arvalid = fetch_io_instRead_arvalid; // @[cpu.scala 98:25]
  assign fetchCrossbar_io_icRead_inst = icache_io_icRead_inst; // @[cpu.scala 137:33]
  assign fetchCrossbar_io_icRead_rvalid = icache_io_icRead_rvalid; // @[cpu.scala 137:33]
  assign fetchCrossbar_io_flashRead_rdata = split64to32_io_data_in_rdata; // @[cpu.scala 138:33]
  assign fetchCrossbar_io_flashRead_rvalid = split64to32_io_data_in_rvalid; // @[cpu.scala 138:33]
  assign split64to32_clock = clock;
  assign split64to32_reset = reset;
  assign split64to32_io_data_in_addr = fetchCrossbar_io_flashRead_addr; // @[cpu.scala 138:33]
  assign split64to32_io_data_in_dc_mode = fetchCrossbar_io_flashRead_dc_mode; // @[cpu.scala 138:33]
  assign split64to32_io_data_out_rdata = flash2Axi_io_dataIO_rdata; // @[cpu.scala 139:33]
  assign split64to32_io_data_out_rvalid = flash2Axi_io_dataIO_rvalid; // @[cpu.scala 139:33]
  assign split64to32_io_data_out_ready = flash2Axi_io_dataIO_ready; // @[cpu.scala 139:33]
  assign memCrossbar_clock = clock;
  assign memCrossbar_reset = reset;
  assign memCrossbar_io_dataRW_addr = memory_io_dataRW_addr; // @[cpu.scala 123:25]
  assign memCrossbar_io_dataRW_wdata = memory_io_dataRW_wdata; // @[cpu.scala 123:25]
  assign memCrossbar_io_dataRW_dc_mode = memory_io_dataRW_dc_mode; // @[cpu.scala 123:25]
  assign memCrossbar_io_dataRW_amo = memory_io_dataRW_amo; // @[cpu.scala 123:25]
  assign memCrossbar_io_mmio_rdata = mem2Axi_io_dataIO_rdata; // @[cpu.scala 141:33]
  assign memCrossbar_io_mmio_rvalid = mem2Axi_io_dataIO_rvalid; // @[cpu.scala 141:33]
  assign memCrossbar_io_mmio_ready = mem2Axi_io_dataIO_ready; // @[cpu.scala 141:33]
  assign memCrossbar_io_dcRW_rdata = dcSelector_io_mem2dc_rdata; // @[cpu.scala 140:33]
  assign memCrossbar_io_dcRW_rvalid = dcSelector_io_mem2dc_rvalid; // @[cpu.scala 140:33]
  assign memCrossbar_io_dcRW_ready = dcSelector_io_mem2dc_ready; // @[cpu.scala 140:33]
  assign memCrossbar_io_clintIO_rdata = clint_io_rw_rdata; // @[cpu.scala 142:33]
  assign memCrossbar_io_plicIO_rdata = plic_io_rw_rdata; // @[cpu.scala 158:25]
  assign tlb_if_clock = clock;
  assign tlb_if_reset = reset;
  assign tlb_if_io_va2pa_vaddr = fetch_io_va2pa_vaddr; // @[cpu.scala 99:25]
  assign tlb_if_io_va2pa_vvalid = fetch_io_va2pa_vvalid; // @[cpu.scala 99:25]
  assign tlb_if_io_mmuState_priv = csrs_io_mmuState_priv; // @[cpu.scala 145:33]
  assign tlb_if_io_mmuState_mstatus = csrs_io_mmuState_mstatus; // @[cpu.scala 145:33]
  assign tlb_if_io_mmuState_satp = csrs_io_mmuState_satp; // @[cpu.scala 145:33]
  assign tlb_if_io_flush = writeback_io_flush_tlb; // @[cpu.scala 134:25]
  assign tlb_if_io_dcacheRW_rdata = dcSelector_io_tlb_if2dc_rdata; // @[cpu.scala 144:33]
  assign tlb_if_io_dcacheRW_rvalid = dcSelector_io_tlb_if2dc_rvalid; // @[cpu.scala 144:33]
  assign tlb_if_io_dcacheRW_ready = dcSelector_io_tlb_if2dc_ready; // @[cpu.scala 144:33]
  assign tlb_mem_clock = clock;
  assign tlb_mem_reset = reset;
  assign tlb_mem_io_va2pa_vaddr = memory_io_va2pa_vaddr; // @[cpu.scala 124:25]
  assign tlb_mem_io_va2pa_vvalid = memory_io_va2pa_vvalid; // @[cpu.scala 124:25]
  assign tlb_mem_io_va2pa_m_type = memory_io_va2pa_m_type; // @[cpu.scala 124:25]
  assign tlb_mem_io_mmuState_priv = csrs_io_mmuState_priv; // @[cpu.scala 147:33]
  assign tlb_mem_io_mmuState_mstatus = csrs_io_mmuState_mstatus; // @[cpu.scala 147:33]
  assign tlb_mem_io_mmuState_satp = csrs_io_mmuState_satp; // @[cpu.scala 147:33]
  assign tlb_mem_io_flush = writeback_io_flush_tlb; // @[cpu.scala 135:25]
  assign tlb_mem_io_dcacheRW_rdata = dcSelector_io_tlb_mem2dc_rdata; // @[cpu.scala 146:33]
  assign tlb_mem_io_dcacheRW_rvalid = dcSelector_io_tlb_mem2dc_rvalid; // @[cpu.scala 146:33]
  assign tlb_mem_io_dcacheRW_ready = dcSelector_io_tlb_mem2dc_ready; // @[cpu.scala 146:33]
  assign dcSelector_clock = clock;
  assign dcSelector_reset = reset;
  assign dcSelector_io_tlb_if2dc_addr = tlb_if_io_dcacheRW_addr; // @[cpu.scala 144:33]
  assign dcSelector_io_tlb_if2dc_wdata = tlb_if_io_dcacheRW_wdata; // @[cpu.scala 144:33]
  assign dcSelector_io_tlb_if2dc_dc_mode = tlb_if_io_dcacheRW_dc_mode; // @[cpu.scala 144:33]
  assign dcSelector_io_tlb_mem2dc_addr = tlb_mem_io_dcacheRW_addr; // @[cpu.scala 146:33]
  assign dcSelector_io_tlb_mem2dc_wdata = tlb_mem_io_dcacheRW_wdata; // @[cpu.scala 146:33]
  assign dcSelector_io_tlb_mem2dc_dc_mode = tlb_mem_io_dcacheRW_dc_mode; // @[cpu.scala 146:33]
  assign dcSelector_io_mem2dc_addr = memCrossbar_io_dcRW_addr; // @[cpu.scala 140:33]
  assign dcSelector_io_mem2dc_wdata = memCrossbar_io_dcRW_wdata; // @[cpu.scala 140:33]
  assign dcSelector_io_mem2dc_dc_mode = memCrossbar_io_dcRW_dc_mode; // @[cpu.scala 140:33]
  assign dcSelector_io_mem2dc_amo = memCrossbar_io_dcRW_amo; // @[cpu.scala 140:33]
  assign dcSelector_io_dma2dc_addr = dmaBridge_io_dcRW_addr; // @[cpu.scala 161:23]
  assign dcSelector_io_dma2dc_wdata = dmaBridge_io_dcRW_wdata; // @[cpu.scala 161:23]
  assign dcSelector_io_dma2dc_dc_mode = dmaBridge_io_dcRW_dc_mode; // @[cpu.scala 161:23]
  assign dcSelector_io_select_rdata = dcache_io_dcRW_rdata; // @[cpu.scala 143:33]
  assign dcSelector_io_select_rvalid = dcache_io_dcRW_rvalid; // @[cpu.scala 143:33]
  assign dcSelector_io_select_ready = dcache_io_dcRW_ready; // @[cpu.scala 143:33]
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io_rw_addr = memCrossbar_io_clintIO_addr; // @[cpu.scala 142:33]
  assign clint_io_rw_wdata = memCrossbar_io_clintIO_wdata; // @[cpu.scala 142:33]
  assign clint_io_rw_wvalid = memCrossbar_io_clintIO_wvalid; // @[cpu.scala 142:33]
  assign plic_clock = clock;
  assign plic_reset = reset;
  assign plic_io_intr_in1 = io_interrupt; // @[cpu.scala 155:25]
  assign plic_io_rw_addr = memCrossbar_io_plicIO_addr; // @[cpu.scala 158:25]
  assign plic_io_rw_wdata = memCrossbar_io_plicIO_wdata; // @[cpu.scala 158:25]
  assign plic_io_rw_wvalid = memCrossbar_io_plicIO_wvalid; // @[cpu.scala 158:25]
  assign plic_io_rw_arvalid = memCrossbar_io_plicIO_arvalid; // @[cpu.scala 158:25]
  assign dmaBridge_clock = clock;
  assign dmaBridge_reset = reset;
  assign dmaBridge_io_dmaAxi_awvalid = io_slave_awvalid; // @[cpu.scala 160:14]
  assign dmaBridge_io_dmaAxi_awaddr = io_slave_awaddr; // @[cpu.scala 160:14]
  assign dmaBridge_io_dmaAxi_awid = io_slave_awid; // @[cpu.scala 160:14]
  assign dmaBridge_io_dmaAxi_awlen = io_slave_awlen; // @[cpu.scala 160:14]
  assign dmaBridge_io_dmaAxi_awsize = io_slave_awsize; // @[cpu.scala 160:14]
  assign dmaBridge_io_dmaAxi_wvalid = io_slave_wvalid; // @[cpu.scala 160:14]
  assign dmaBridge_io_dmaAxi_wdata = io_slave_wdata; // @[cpu.scala 160:14]
  assign dmaBridge_io_dmaAxi_wstrb = io_slave_wstrb; // @[cpu.scala 160:14]
  assign dmaBridge_io_dmaAxi_bready = io_slave_bready; // @[cpu.scala 160:14]
  assign dmaBridge_io_dmaAxi_arvalid = io_slave_arvalid; // @[cpu.scala 160:14]
  assign dmaBridge_io_dmaAxi_araddr = io_slave_araddr; // @[cpu.scala 160:14]
  assign dmaBridge_io_dmaAxi_arid = io_slave_arid; // @[cpu.scala 160:14]
  assign dmaBridge_io_dmaAxi_arlen = io_slave_arlen; // @[cpu.scala 160:14]
  assign dmaBridge_io_dmaAxi_arsize = io_slave_arsize; // @[cpu.scala 160:14]
  assign dmaBridge_io_dmaAxi_rready = io_slave_rready; // @[cpu.scala 160:14]
  assign dmaBridge_io_dcRW_rdata = dcSelector_io_dma2dc_rdata; // @[cpu.scala 161:23]
  assign dmaBridge_io_dcRW_rvalid = dcSelector_io_dma2dc_rvalid; // @[cpu.scala 161:23]
  assign dmaBridge_io_dcRW_ready = dcSelector_io_dma2dc_ready; // @[cpu.scala 161:23]
endmodule
